MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �N��u ��u ��u �O;���u ڳ���u ڳ�ڰu �����u ��u!ږu ڳ���u ڳ���u ڳ���u �Rich�u �                        PE  L �=�L        � !
  :  v      ��     P                           ��                      �� M   ā (    � �                   � x                                  @w @            P                           .text   8     :                   `.rdata  �7   P  8   >             @  @.data   D2   �     v             @  �.rsrc   �   �     �             @  @.reloc  �'   �  (   �             @  B                                                                                                                                                                                                                                                                                                                                                U����V��H�QV�ҡ���U�H�E�IRj�PV�у���^]� ���������̡���P�BQ��Y�U��j�h�Ed�    P���8�3�P�E�d�    �F   ��uh����H�A�U�R�Ћ���Q�Jj j��E�hPQP�эU�R�E�    ��&  ����H�A�U�R�E������Ѓ�3��M�d�    Y��]ø   �M�d�    Y��]�����������������������U��E�� tHt3�]ùģ�4J  �����]ø   ]������U��V������M�$�jn �F�$�]�\n �}���m ^]� ������������U�����E�P�E���   ���$P��]� ������������U�����E�P�E�R,���$P��]� ���������������U�������   ���   ]����������̡���P@�B,Q�Ѓ����������������U�����PH�EP�EPQ���   �у�]� �������������U�����PH�EPQ���   �у�]� ̡���PH���   h�  Q�Ѓ�������̡���PH���   j h�  Q�Ѓ�����̡���PH���   h�  Q�Ѓ�������̡��V��Hl�V�AR�Ѓ��F    ^�U��j�h�Ed�    P��4SV�8�3�P�E�d�    3�;���  �]��]ĉ]ȉ]̉]Љ]؉]ԡ�����   �Sj�]��Ћ���Q�J���E�P�ы���B�PSj��M�h�QQ�҃�������   �R|�E�P���E��ҡ���H�A�U�R�]��������U��U���]�E܋QH�RP���������U��U���]�PH�R �E�P�ҋE�M�Qh�   �uĉE��%  ����tk�U�R�s  ������   �M؋��   ��S�Ћ���Eċ��   ���   �E�P�ы�����   ���   �M�Q�ҍE�Ph�   �$  ����u^������   ���   �E�P�ы�����   ���   �M�Q�ҍE�P��r  ���M��E������B:  3��M�d�    Y^[��]Ë�����   �M؋��   S�ЍM�Q���r  ������   ���   �M�Q�ҡ�����   ���   �U�R�Ѓ��M��E�������9  �ƋM�d�    Y^[��]���������U�����UVW���H@�A,R�Ћ���Q���B ������=ݣ �g  �����Q�B,���$h�  ���Ћ���Q�B4jh�  ������Q����Q�B,���$h�  ���Ћ���Q�B0j h�  ���Ћ���Q�B4j h�  ���Ћ���Q�B4j h�  ���������Q�B,���$h�  �����xQ��Q����Q�B,�5pQ�����$h�  �������Q�B,���$h�  ���������Q���$h�  �B,���Ћ���Q�B0jh�  ���������Q�B,���$h�B ���Ћ���Q�B$hݣ �����G    �G    _�   ^]� ��������U�����H@�U�A,VWR�Ћ���Q��j �ȋ��   h�  �Ћuj �΋��?L  �8�  u��t��u_3�^]� j ���L  �8�  u��u�_�   ^]� �����U��S�ًMhݣ ��M  ��tBV�u�����H@�Q,W�}W�ҡ�����   �BT�����ЋMVQW���N�  _^[]� 3�[]� U��j�hFd�    P��pSVW�8�3�P�E�d�    �M܋u3�;���  ����HH���   h�  V�҃�����  j�}�}�I�  ���E��}�;�t���h  �؉]���}�ߡ���HH���   h�  V�E������ҋ�����HH���   j h�  V�҉E����HH���   h�  V�ҋM���R��j WQP���ҡ���HH���   h�  3�V�}��҃�����  �}����Hl�UR�S�E�P�AWR����E���Uă����U����U��������؅��c  �E�    �
���������؋M�U��<�����HH���   j h�  V�����L�T���G�EС��j �MԋHH�U؋��   h�  V�ҋMЋ���I�<ȋBH���   j h�  V�ыM؍I�Ѝ��'j h�  V�]��@�g�]��@����g�HH���   �]��ҋ���[�<ȋBH���   j h�  V�ыMԍI�Ѝ��'��<�@�g�@�g���E������E��������U��E������������U��������������U��������������������c ��������������Dz
��������������E����E����E������������E��E�@�E��U����E��U����E��U�;E�c����}��ʋ]����E����������D{���������U��������U��������U�������������U����U����U�����������������������b ��������������Dz��������������E������M����M����ʋM��ʋQ�E���Q���\�I�\��E������E�BH���   h�  GV�}��у�;��-�������Bl�K�PQ�҃��C    �M�d�    Y_^[��]� ���������U��Q�E�M���������D��   �y ��   ����HH���   S�]VWj h�  S�ҋ����HH���   h�  S3��҃���~_3���E��F�@�Fh�  �E����G����D����D��E��P�����������^��^��^�����QH���   �у�;�|�_^[��]� �������+E  �����������V��V觍  ���    ^�������������U��j�hYFd�    PQV�8�3�P�E�d�    �E�    ����H�u�QV�E�    �ҡ���H�U�AVR�Ѓ�����Q�B<���E�    �E�   �Ћ���Q�M�RLj�j�QP���ҋƋM�d�    Y^��]����������������U��V���5~  �Et	V�Ɇ  ����^]� ���������������U��j�h�Fd�    P��t  SVW�8�3�P�E�d�    �M̋}3�;���  ������   �BT���Ћ���Q@���B,W�Ћ���Q��SV�ȋBlh�  �Ћ��u�;��r  ������   �Bt���Ѕ��W  ������   �B4���ЉE�;��  h  ��h  �����}�;��  ������   �Bt���Ћ���Q@�EԋB,W�Ћ���Q�MԋRp��Qh�  ����ShTR�M������������   �Bt�Ή]��Ћ�����   �ȋBx�ЍM�QP�U�R�������������   P�B|���E��Ћ���Q�J�E�P�]��ы���B�P�M�Q�E������ҡ�����   �E�RD��P���ҡ�����   �Bt���Ћ���QH�R,������Q���ҋ����   �������PH�u�R0������P���ҡ�����   �BSj���Љ�p�����t�����x�����|����]��]��]��M��E�   �A  �]��]��E��<�  �E�h  �E��]܉]��]�]ȉ]ԉ]�3��g  ���E�;���  ������   �M�BT�Ћ��}�;��  ��聜  ��u���ŋ  ;E�u	�U�R��  ������   �}��Bt����ShE  ���5���;�tW�����Q@P�B,�Ћ���Q���ȋB$V�Ћ�����   �Bt��F�Ћ���QHVhE  P���   �Ѓ�;�u�������   �Bt����j��������E�;���   ������   �Bt���Ћ�����   �ȋB4�Ћ�;���   �I 9]���   ������   �B����=%  tb=+F t[=  tT=�  tM=  tF=  t?=  t8=  t1=	  t*=  t#=  t=  t=  t=  t=%G u����QH���   jV�Ѓ��E؋�����   �B(���Ћ�;��D����u��M�Q�����  � �]����@�]��4�  �E��Eȃ��M��$�����u�E��Eȃ����]����$h�B �P�����������E�����������D{"���$h�B ���E�   � ������������؋E�MSS�U�RjPQ���k  �E�;��0  9]�u|9]�t�U�R耵  ��9]�t�E�P诬  ������Q@�EЋJP�эU�R�E��M�  ���M��]��E��>  ��p����E������+  �EȋM�d�    Y_^[��]� ���k�����;�u	�E�P�  ����Q���   Sh�  ���Ћ�;�}3��
��~�   ����Q�B4Wh�  ���ЋM�Q�M��������ShLR�M��E������������   �P|�M�Q�M��E��ҡ���H�A�U�R�E��ЋM����  ������   �M�P�BD�Ѝ�@������  ����Q�B0jh2  ��@����E��Ћ���Q�B4Wh5  ��@����Љ�`�����d�����l�����h����M�E艍T�����T���Q��@���h�   �E���\�����X����)  ����u#��T����E��*  ��@����E�贮  �,	  ��l���R�������h���P�����Ẻx��P�E�%|  �M���*���3ɋ��   �������Q�B~  ��;�t�W�;�|��H�Q��J�Q��Q�y����3��M�����B�P��@����ҍ�T����E��R)  ��@����E���  9]��w  j��|  ���E�E�;�t���[  �E��]�Ë}�Eԋ ��S���E��E�����P������P���Z����MP�E���ҋESP���3j  �ωE��iQ  ���r�  h�  �M��I  P�M��E�	�x=  �M��E��;  �M���������Q�ȋB ��PhE  �������E�;�t������   �R�M�Qj���ҋM̋���   W��h�  ��`  ����;��o  ����$��h�  �������$h�  ����������������$h�  ���q������$h�  �����������������$h�  ���D������$h�  ���������[�������$h�  ���������$h�  ���������.�������P���   Sh�  ���Ћϋ��]�������QS�ȋB0h�  �Ћ���Q���   j h�  ���Ћϋ��$�������QS�ȋB4h�  �Ћ���Q���   j h�  ���Ћϋ����������QS�ȋB4h�  �Ћ���Q���   j h�  ���Ћϋ���������QS�ȋB4h�  �Ћ���Q���   j h�  ���Ћϋ��y�������QS�ȋB4h�  �Ћ���Q���   j h�  ���Ћϋ��@�������QS�ȋB4h�  �Ћ���Q���   j h�  ���Ћ؋���������QS�ȋB4h�  �Ћ���Q���   j h�  ���ЉE��E������$h�  �������h�������Q���   j h�  ���ЉE��E������$h�  �������/�������Q���   j h�  ���ЉE��E������$h�  �M��������������Q���   j h�  ���ЉE��E������$h�  ��������������Q���   j h�  ���Ћ؋����������QS�ȋB0h�  �Ћ���Q���   j h�  ���Ћϋ���������QS�ȋB0h�  �Ћ���Q���   j h�  ���Ћϋ��x�������QS�ȋB0h�  �Ћ���Q���   j h�  ���Ћϋ��?�������QS�ȋB0h�  �Ћ�����   �EЋRDP���ҋMj h�  �#����؅���   j h�  ���+K  j h�  ��������E���  �����������Qj �ȋ��   h�  �ЋM�E���������Q�M��R0Qh�  ���ҋ���������Qj �ȋ��   h�  �ЋM�E��a�������Q�M��R0Qh�  ��������$h�  ���4����������M���$h�  ���������������$��h�  �����M̋�]苐�   ���$S�ҋE썍p���Qh�   ��t�����p�����  ������  ������   �P4���ҋ؅���  ������   �BL����j h@R�M�����������   �R|�E�P���E�
�ҡ���H�A�U�R�E��Ћ�����   �M�BL���Ћ���Q���   j h�  ���ЋˉE���������Q�M��R0Qh�  ���ҡ���P���   j h�  ���ЋˉE����������Q�M��R4Qh�  ��������$h�  ���+������$h�  ���������B�������P���   j h�  ���ЋˉE��o�������Q�M��R4Qh�  ���ҡ���P���   j h�  ���Ћˋ��4�������QV�ȋB4h�  �Ћ�����   �Bj j���Ћ�����   �BDW���Ћ�����   �Bj j����h  �bY  ��������   3�9]�t�M�Q�U�  ��9]�t�U�R脡  ���E�;�t����Q@P�B�Ѓ��M�;�t�L����E�;�t����Q@P�B�Ѓ��E�;�t����Q@P�B�Ѓ��M�Q�E���{  ���M��]��E��;3  ��p����E������   3��M�d�    Y_^[��]� ������   �M�PT�ҋM�����������Qj S�ȋBlh�  �Ћ΋����������QS�ȋBph�  ��j h0R�M�����������   �R|�E�P���E��ҡ���H�A�U�R�E��Ѓ�j���#E  ������   �BDW���Ѓ}� t�M�Q��  ���}� t�U�R��  ������H@�U�AR�ЋM�����������Q@�EȋJP�эU�R�E��z  ���M��E�    �E���1  ��p����E�������  �EЋM�d�    Y_^[��]� �U��j�h)Gd�    PQV�8�3�P�E�d�    h`Rjh�j��t  �����u�3��E�;�t���Qk  ��Q�ƋM�d�    Y^��]����������U��j�hpGd�    P��4V�8�3�P�E�d�    ����H�A�U�R�Ћ���Q�Jj j��E�h�RP�у�����B�P<�M��E�    �҅�u0����H�A�U�R�E������Ѓ��   �M�d�    Y^��]Ë���Q�J�E�P�ы���B�Pj j��M�h�RQ�ҡ���H�A�U�R�E��Ћ���Q�Jj j��E�h�RP�у�(�U�R�M��E��l  � j P�E�PhP0 j�M�Qhݣ �E��}�  ���M����E��m  ����B�P�M�Q�E��ҡ���H�A�U�R�E� �Ћ���Q�J�E�P�E������у��ƋM�d�    Y^��]����U��E���� ]��U�����P8�EPQ�JD�у�]� ���̡���H8�Q<�����U�����H8�A@V�u�R�Ѓ��    ^]�������������̡���H8�������U�����H8�AV�u�R�Ѓ��    ^]��������������U�����P8�EP�EP�EPQ�J�у�]� ������������U�����P8�EP�EPQ�J�у�]� ����P8�BQ�Ѓ����������������U�����P8�EPQ�J �у�]� ����U�����P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U�����P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�����P8�EP�EPQ�J(�у�]� U�����P8�EP�EP�EPQ�J,�у�]� ������������U�����P8�EP�EP�EPQ�J�у�]� ������������U�����P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�����P8�EP�EPQ�J0�у�]� U�����P8�EP�EP�EPQ�J4�у�]� ������������U�����P8�EPQ�J8�у�]� ����U�����H��x  ]��������������U�����H��|  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H�A,]�����������������U�����H�QV�uV�ҡ���H�Q8V�҃���^]�����̡���H�Q<�����U�����H�I@]����������������̡���H�QD����̡���H�QH�����U�����H�AL]�����������������U�����H�IP]�����������������U�����H��<  ]��������������U�����H��,  ]��������������U�����H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡���H���   �����H���  ��U�����H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U�����H�A]�����������������U�����H��\  ]��������������U�����H�AT]�����������������U�����H�AX]�����������������U�����H�A\]����������������̡���H�Q`����̡���H�Qd����̡���H�Qh�����U�����H�Al]�����������������U�����H�Ap]�����������������U�����H�At]�����������������U�����H��D  ]��������������U�����H��  ]��������������U�����H�Ix]�����������������U�����H��@  ]��������������U��V�u����  ����H�U�A|VR�Ѓ���^]���������U�����H���   ]��������������U�����H��h  ]��������������U�����H��d  ]��������������U�����H���  ]�������������̡���H���   ��U�����H��l  ]��������������U�����H��   ]��������������U�����H��  ]��������������U��V�u����  ����H���   V�҃���^]���������̡���H��`  ��U�����H��  ]��������������U�����H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U�����H���  ]��������������U��U�E����H�E���   R���\$�E�$P�у�]�U�����H���   ]��������������U�����H���   ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���   ]��������������U�����H���   ]��������������U�����H���   ]��������������U�����H���   ]��������������U�����H���   ]��������������U�����H���   ]��������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�����H��8  ]��������������U��V�u(V�u$�E�@����R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@����R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�����P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�����P0�EP�EP�EP�EPQ���   �у�]� ����̡���P0���   Q�Ѓ�������������U�����P0�EP�EPQ���   �у�]� �������������U�����P0�EP�EP�EP�EPQ���   �у�]� ����̡���P0���   Q�Ѓ������������̡���H0���   ��U�����H0���   V�u�R�Ѓ��    ^]�����������U�����H��H  ]��������������U�����H��T  ]�������������̡���H��p  �����H���  ��U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ������   �Qj PV�ҡ�����   ��U�R�Ѓ� ��^��]��������U���4VhLGOg�M��|�  ����Q��X  3�VP�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�у� �M��b�  ������   �PT�M�Q�҃���u'�u���ܑ  ������   ��U�R�Ѓ���^��]Ë�����   �JT�E�P�ыu��P���ܑ  ������   ��M�Q�҃���^��]���������������U�����H��  ]��������������U�����H��\  ]��������������U�����H�U��t  ��V�uVR�E�P�у���胜  �M�軛  ��^��]�����U�����H�U���  ��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]����������������U�����H�U���  ��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]����������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H�U�E��VWj R�UP�ERP��t  �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�(_��^��]��U�����H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у�$��^��]���U�����H��8  ]��������������U���  �8�3ŉE��M�EPQ������h   R�{ ����x	=�  |#�����H��0  h�RhF  �҃��E� ����H��4  ������RhS�ЋM�3̓��C8 ��]�������U�����H��  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]����U�����H��  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]����U�����H��p  ��4�҅���   h���M���  ����P�E�R4Ph���M��ҡ���P�E�R4Ph���M��ҡ���H��X  j �U�R�E�hicMCP�ы���E�    �E�    ���   j P�A�U�R�Ћ�����   �
�E�P�ы�����   ��M�Q�҃�$�M�諌  ��]��������U�����H��p  ��4V�҅�u����H�u�QV�҃���^��]�Wh!���M���  ����P�E�R4Ph!���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �PH�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ�����   ��U�R�Ѓ�4�M�蝋  _��^��]������U�����H��p  ��4V�҅�u����H�u�QV�҃���^��]�Wh����M���  ����P�E�R4Ph����M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �PH�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ�����   ��U�R�Ѓ�4�M�荊  _��^��]������U�����H��p  ��4�҅�u��]�Vh#���M���  ����P�E�R4Ph#���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �P8�M�Q�ҋ������   ��U�R�Ѓ�(�M�赉  ��^��]���������������U�����H��p  ��4�҅�u��]�Vhs���M��4�  ����P�E�R4Phs���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �P8�M�Q�ҋ������   ��U�R�Ѓ�(�M��Ո  ��^��]���������������U�����H���  ]��������������U�����H��@  ]��������������U�����H���  ]��������������U��V�u���t����QP��D  �Ѓ��    ^]������U�����H��H  ]��������������U�����H��L  ]��������������U�����H��P  ]��������������U�����H��T  ]��������������U�����H��X  ]��������������U�����H��\  ]�������������̡���H��d  ��U�����H��h  ]��������������U�����H��l  ]�������������̡���H���  ��U�����H�U���  ��VR�E�P�ыu��P���Æ  �M��ۆ  ��^��]�����U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H���  ]��������������U�����H��$  ]��������������U�����H��(  ]��������������U�����H��,  ]�������������̡���H��0  �����H��<  ��U�����H���  ]�������������̡���H���  ��U�����H���  ]������������������������������U�����H��  ]�������������̡���H��P  �������   ���   ��Q��Y��������U�����H�A�U��� R�Ћ���Q�Jj j��E�hSP�ы���B�P�M�Q�ҡ���H�I�U�R�E�P�ы���B�P<�� �M��ҋ���Q�M�RLj�j�QP�M��ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�҃���]��������������U��E��u�ģ�MP�EPQ�  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3hSj;h�j�U  ����t
W���~�  �3��F��u_^]� �~ t3�9_��^]� ����H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ����H<�Q��3Ʌ����^��������������̃y t�   ËA��uË���R<P��JP�у��������U����u����H�]� ����J<�URP�A�Ѓ�]� ���������������U��ģ��u����H�]Ë���J<�URP�A�Ѓ�]�U��ģ��$V��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�SP�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���[t.����B�u�HV�ы���B�P�M�Q�҃���^��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^��]���������������U��ģ��$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]����������������U��ģ��$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]��U��ģ��$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�hHSP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]����U�����H<�A]����������������̡���H<�Q�����V��~ u>���t����Q<P�B�Ѓ��    W�~��t���ڂ  W�TI  ���F    _^��������U���V�E�P��讔  ��P�������M��虂  ��^��]��̃=̣ uK�ģ��t����Q<P�B�Ѓ��ģ    �У��tV���P�  V��H  ���У    ^������������U���H����H�AS�U�V3�R�]��Ћ���Q�JSj��E�hLSP�ы���B<�P�M�Q�ҋ����H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��8�  �M�Q�U�R�M�舠  ���&  W�}�}���   ������   �U��ATR�Ћ�������   ����Q�J�E�P���ы���B���   ���M�Qj�U�R���Ћ���Q�J���E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Bx��W�M����E���t�E� ��t����Q�J�E�P����у���t����B�P�M�Q����҃��}� u"�E�P�M�Q�M��s�  ��������E�_^[��]ËU��U�_�E�^[��]��U���DSV�u3ۉ]�;�u_����H�A�U�R�Ћ���Q�JSj��E�hLSP�ы���B<�P�M�Q�ҋ����H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��q�  �M�Q�U�R�M����  ���p  W�}��I �E����   ������   �U��ATR�Ћ�������   ����Q�J�E�P���ы���B���   ���M�Qj�U�R���Ћ���Q�J���E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Bx��W�M����E��t�E ��t����Q�J�E�P����у���t����B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*������   P�BH�Ћ���Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��b�  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��Ü  �EP�M�Q�M�u��u��  ����   �u���E���tA��t<��uZ������   �M�PHQ�ҋ���Q���ȋBxV�Ѕ�u-�   ^��]Ë�����   �E�JTP��VP�[�������uӍUR�E�P�M�脜  ��u�3�^��]����������V��~ u>���t����Q<P�B�Ѓ��    W�~��t���Z}  W��C  ���F    _^��������hԣPhD 萜  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��hԣjhD 輛  ����t
�@��t]��3�]��������Vhԣj\hD ��茛  ����t�@\��tV�Ѓ���^�����Vhԣj`hD ���\�  ����t�@`��tV�Ѓ�^�������U��VhԣjdhD ���)�  ����t�@d��t
�MQV�Ѓ�^]� ������������U��VhԣjhhD ����  ����t�@h��t
�MQV�Ѓ�^]� ������������VhԣjlhD ��謚  ����t�@l��tV�Ѓ�^�������U��Vhԣh�   hD ���v�  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vhԣh�   hD ���&�  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhԣjphD ���ٙ  ����t�@p��t�MQV�Ѓ�^]� �أ^]� ��U��VhԣjxhD ��虙  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��VhԣjxhD ���Y�  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��VhԣjxhD ����  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������hԣjhD 还  ����t	�@��t��3��������������U��V�u�> t+hԣjhD 胘  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0hԣjhD �A�  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��VhԣjhD �����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��VhԣjhD ��蹗  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vhԣj hD ���|�  ����t�@ ��tV�Ѓ�^�3�^���Vhԣj$hD ���L�  ����t�@$��tV�Ѓ�^�3�^���U��Vhԣj(hD ����  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vhԣj,hD ���ɖ  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vhԣj(hD ��艖  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vhԣj4hD ���<�  ����t�@4��tV�Ѓ�^�3�^���U��Vhԣj8hD ���	�  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vhԣj<hD ��蹕  ����t�@<��t
�MQV�Ѓ�^]� ������������VhԣjDhD ���|�  ����t�@D��tV�Ѓ�^�3�^���U��VhԣjHhD ���I�  ����t�M�PHQV�҃�^]� U��VhԣjLhD ����  ����u^]� �M�PLQV�҃�^]� �����������U��VhԣjPhD ���ٔ  ����u^]� �M�U�@PQRV�Ѓ�^]� �������VhԣjThD ��蜔  ����u^Ë@TV�Ѓ�^���������U��VhԣjXhD ���i�  ����t�M�PXQV�҃�^]� U��Vhԣh�   hD ���6�  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vhԣh�   hD ����  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vhԣh�   hD ��薓  ����u^]� �M���   QV�҃�^]� �����U��Vhԣh�   hD ���V�  ����u^]� �M���   QV�҃�^]� �����U��Vhԣh�   hD ����  ����u^]� �M���   QV�҃�^]� �����U��Vhԣh�   hD ���֒  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vhԣh�   hD 蕒  ����u����H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]��U��Vhԣh�   hD ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vhԣh�   hD ��趑  ����t���   ��t�MQ����^]� 3�^]� �U��Vhԣh�   hD ���v�  ����t���   ��t�MQ����^]� 3�^]� �U��Vhԣh�   hD ���6�  ����t���   ��t�MQ����^]� 3�^]� �Vhԣh�   hD �����  ����t���   ��t��^��3�^����������������U��Vhԣh�   hD ��趐  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vhԣh�   hD ���f�  ����t���   ��t�MQ����^]� ��������U��Vhԣh�   hD ���&�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vhԣh�   hD ���ُ  ����t���   ��t��^��3�^����������������VW��3����$    �hԣjphD 菏  ����t�@p��t	VW�Ѓ���أ�8 tF��_��^�������U��SW��3�V��    hԣjphD �?�  ����t�@p��t	WS�Ѓ���أ�8 tqhԣjphD ��  ����t�@p��t�MWQ�Ѓ�����أhԣjphD �ێ  ����t�@p��t	WS�Ѓ���أV���7�����tG�]����E^��t�8��~=hԣjphD 莎  ����t�@p��t	WS�Ѓ���أ�8 u_�   []� _3�[]� ����������U��Vhԣj\hD ���9�  ����t3�@\��t,V��hԣjxhD ��  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vhԣj\hD ���ٍ  ����t3�@\��t,V��hԣjdhD 跍  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vhԣj\hD ���v�  ����tG�@\��t@V�ЋEhԣjdhD �E��E�    �E�    �@�  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vhԣj\hD �����  ����t\�@\��tUV��hԣjdhD �׌  ����t�@d��t
�MQV�Ѓ�hԣjhhD 讌  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vhԣj\hD ���i�  ������   �@\��t~V��hԣjdhD �C�  ����t�@d��t
�MQV�Ѓ�hԣjhhD ��  ����t�@h��t
�URV�Ѓ�hԣjhhD ��  ����t�@h��t
�MQV�Ѓ���^]� ��U���VhԣjthD ��趋  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���hԣj`hD �~�  ����th�@`��ta�M�Q�Ѓ���^��]� hԣj\hD �M�  �u����t4�@\��t-V��hԣjdhD �(�  ����t�@d��thأV�Ѓ���^��]� ������U���Vhԣh�   hD ����  ����tR���   ��tH�MQ�U�R���ЋuP���k���hԣj`hD 誊  ����t|�@`��tu�M�Q�Ѓ���^��]� hԣj\hD �E�    �E�    �E�    �d�  �u����t3�@\��t,V��hԣjdhD �?�  ����t�@d��t
�U�RV�Ѓ���^��]� ��������������U�����E�PH�B���$Q�Ѓ�]� ���������������U�����PH�EPQ���   �у�]� �U�����PH�EPQ���  �у�]� �U�����PH�EPQ���  �у�]� �U�����PH�EP�EPQ��  �у�]� �������������U�����PH�EP�EPQ��  �у�]� ������������̡���PH���  Q�Ѓ�������������U�����PH�EPQ���  �у�]� ̡���PH���   j Q�Ѓ�����������U�����PH�EPj Q���   �у�]� ��������������̡���PH���   jQ�Ѓ�����������U�����PH�EPjQ���   �у�]� ��������������̡���PH���   jQ�Ѓ����������U�����PH�EPjQ���   �у�]� ���������������U�����PH�EP�EPQ���   �у�]� �������������U�����PH�EP�EPQ���   �у�]� ������������̡���PH���   Q�Ѓ�������������U�����PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���a  ������t�E����QH���   PVW�у���_^]� �����U��EVW���MPQ�a  ������t�M����BH���   QVW�҃���_^]� ̡���PH���   Q�Ѓ������������̡���PH���   Q�Ѓ�������������U�����PH�EPQ���   �у�]� �U�����PH�EPQ���   �у�]� �U�����PH�EP�EPQ��8  �у�]� �������������U�����PH�EP�EPQ��   �у�]� ������������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ������������̡���PH��  Q�Ѓ������������̡���PH��  Q�Ѓ�������������U�����PH�EP�EPQ��  �у�]� �������������U�����PH�EP�EP�EPQ��   �у�]� ���������U�����PH�EP�EP�EP�EPQ��|  �у�]� �����U�����PH�EPQ��  �у�]� ̡���PH��T  Q�Ѓ�������������U�����PH�EP�EPQ��  �у�]� �������������U�����PH�EPQ��8  �у�]� �U�����PH�EPQ��<  �у�]� �U�����PH�EPQ��@  �у�]� �U�����PH�EP�EP�EPQ��D  �у�]� ��������̡���PH��L  Q��Y��������������U�����PH�EPQ��H  �у�]� ̡��V��H@�Q,WV�ҋ���Q��j �ȋ��   h�  �Ћ���QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡���P@�B,Q�Ћ���Q��j �ȋ��   h�  �������U�����E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�����E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�����PH�EP�EP�EPQ��   �у�]� ��������̡���HH��  ��U�����HH��  ]��������������U�����E�PH��$  ���$Q�Ѓ�]� �����������̡���PH��(  Q�Ѓ�������������U�����PH�EP�EPQ��,  �у�]� �������������U�����E�PH�EP�E���$PQ��0  �у�]� ���̡���PH���  Q�Ѓ������������̡���PH��4  Q�Ѓ������������̋��     �������̡���PH���|  jP�у���������U�����UV��HH��x  R��3Ƀ������^��]� ��̡���PH���|  j P�у��������̡���PH��P  Q�Ѓ������������̡���PH��T  Q�Ѓ������������̡���PH��X  Q�Ѓ�������������U�����PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡���PH��`  Q�Ѓ�������������U�����PH�EPQ��d  �у�]� �U�����E�PH��h  ���$Q�Ѓ�]� ������������U�����E�PH��t  ���$Q�Ѓ�]� ������������U�����E�PH��l  ���$Q�Ѓ�]� ������������U�����PH�EPQ��p  �у�]� �U�����PH�EP�EP�EP�EPQ���  �у�]� �����U�����PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U�����E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E����HH�E���   R�U���$P�ERP�у�]����������������U���E�M�XS�<�  �M;�|�M;�~��]�����������U�����PH�E���   Q�MPQ�҃�]� ������������̡���PH���   Q��Y�������������̡���PH���   Q�Ѓ������������̡���PH���   Q��Y��������������U�����PH�EP�EPQ���   �у�]� �������������U�����PH�EP�EP�EP�EP�EPQ���  �у�]� ̡���PH��t  Q��Y�������������̋�� dS�@    ��dS����Pl�A�JP��Y��������U����V��Hl�V�AR�ЋE����u
�   ^]� ����Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË���QlP�B�Ѓ�������U�����Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E����HH�ER�U���$P���  R�Ѓ�]����U�����HH���  ]��������������U�����HH���  ]��������������U��U0�E(����HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U�����HH���  ]��������������U�����E�PH�EP���$Q���  �у�]� ��������U���SV���L  �؉]����   �} ��   ����HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}���L  ����   �]��I �E�P�M�Q�MW�M  ��t_�u�;u�W�I ������u�E����ҋL�;L�t-����Bl�S�@����QR�ЋD������t	�M�P�eL  F;u�~��}��MG�}��0L  ;��x����]�_^��[��]� ^3�[��]� U������SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u����HH���  �'��u����HH���  ���uš���HH���  S�ҋȃ��E��t�W�L  ����HH���   h�  S3��҃����  ���_�u����    ����Hl�U�B�IWP�ы�������   ����F�J\�UP�A,R�Ѓ���t�K�Q�M�%K  ����F�J\�UP�A,R�Ѓ���t�K�Q�M��J  �E��;Pt&�F����Q\�J,P�EP�у���t	�MS��J  ����v�B\�M�P,VQ�҃���t�M�CP�J  ����QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U�����HH���   ]�������������̡���PH���   Q��Y��������������U�����HH���  ]��������������U������P���   V�uW�}���$V�����E������At���E������z����؋���Q�B,���$V����_^]����������������U���0�����U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١���]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U�����HH�]��U�����H@�AV�u�R�Ѓ��    ^]�������������̡���HH�h�  �҃�������������U�����H@�AV�u�R�Ѓ��    ^]��������������U�����HH�Vh  �ҋ�������   �EPh�  ��O  ����t]����QHj P���   V�ЋMQh(  ��O  ����t3����JH���   j PV�ҡ�����   �B��j j���Ћ�^]á���H@�QV�҃�3�^]�������U�����H@�AV�u�R�Ѓ��    ^]��������������U�����HH�Vh�  �ҋ�����u^]á���HH�U�E��  RPV�у���u����B@�HV�у�3���^]�������U�����H@�AV�u�R�Ѓ��    ^]��������������U�����HH�I]�����������������U�����H@�AV�u�R�Ѓ��    ^]��������������U�����PH�EPQ���  �у�]� �U�����PH�EPQ���  �у�]� ̡���PH���  Q�Ѓ�������������U�����HH���  ]��������������U�����E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡���PH���  Q�Ѓ�������������U�����PH�EP�EPQ���  �у�]� ������������̡���PH��  Q�Ѓ�������������U�����PH�EP�EP�EPQ���  �у�]� ��������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ�������������U�����PH�EPQ��  �у�]� �U�����PH�EPQ��  �у�]� ̋������������������������������̡���HH���  ��U�����HH���  ]��������������U�����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U�����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡���PH��,  Q�Ѓ�������������U�����PH�EPQ��X  �у�]� ̡���PH��\  Q�Ѓ�������������U�����HH��0  ]��������������U������W���HH���   j h�  W�҃��} u�   _��]� Vh�  �oJ  ��������   ����HH���   j VW�҃��M��E  ����P�E�R0Ph�  �M����E����P�B,���$h�  �M��Ћ���Q@�J(j �E�PV�у��M��E  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7����U�HH���   RW�Ѓ���u����QH���   jW�Ѓ���t�   �����   ����QH���   W�Ѓ��} u(����E�QH�M���  P�ESQ�MPQW�҃��B�u��t;����U�HH�ER�USP���  VRW�Ћ�����   �B(�����Ћ���uŃ; u����QH���   W�Ѓ���t3���   �W��u1����QH���   �Ћ���E�QH���   PW�у�_^[]� ����BH���   �у��} u0����M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ����QH�h  �Ћ؃���u_^[]� ������   �u�Bx���Ћ�����   P�B|���Ѕ�tU����E�QH�MP�Ej Q���  VPW�у���t������   �ȋBHS�Ћ�����   �B(���Ћ���u�_^��[]� ��������������U��EV���u����HH���  �'��u����HH���  ���u����HH���  V�҃���u3�^]� P�EP���N���^]� ���������U���D����HH���   S�]VWh�  S�ҋ����HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��>
  ������   �B���Ћ��=�  �  �QH���   Wh:  S�Ћ���QH�E����   h�  S�Ћ���QHW�����   h�  S�uԉ}��Ћ���QH�E苂  S�Ћ���QH�EЋ��  S�Ѓ�(�E��E�pS��~~�M���M�I �MЅ�tMj�W衁  ���t@�@�Ẽ|� �4�~����%�������;�u/��� �  ;E�~�E؋���  E���E�;Pu�E���E��E�G;}�|��}� ��   �u�j S���gE  ����  ���H  ��ti����B  �}�;�u^����H���  �4�htS��h�  V�҃��E���b  �M��E��iH  ��t�}� t��tVP�E�P��  ����}܋���Q���  �4�htS��h�  V�Ѓ��E����  �M�3�;�t;�tVQP���  ���E�;�~-����QhtS��h�  P���   �Ѓ��E�;���  ����E��QH��  j�PS�у�����  �u�;�tjS���5D  ���{  ���G  �E���}����BH���   Wh�  S�у�3��E�}�9}��]  �}���}����$    �MЅ��J  �U�j�R�  ����6  �M̍@�|� ���]�~����%�������9E���  ���͈  �E�3�3ɉE܉M�9C��   ��$    �����������ti�]������������M�ҋ9�<��}�҉T��y�]��|��]��z�|��y�]��|��]��z�|��I�}��]��L��M��}ȃ��T����M�A�M�;K�v����E؅��0  �+U�j��PR�M��l  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t4�U�M��@���P�Q�P�Q�P�Q�P�Q�@�A�M��Eȍ@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A;]�}_�UȋE�9�uT�ȋL�����������w0�$�t� �U���4���M���t���U���t��	�M���t��M���;]�|��E܃�F�M�;]������U�;U��  �U�R�9  �E�P�0  �M�Q�'  ��_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q�P �Q�P$�Q�P(�I�H,��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@���E��}�;E�������U�R�	  �E�P�	  ���  ���   �B����=  ��  ����QH���   j h(  S�Ћ���QH�����   h(  S�ЋЃ�3��U؅�~"��ǅ�t�|� t�4N��tN�@;�|�u��u܋���Q���  �4v�htS��hK  V�Ѓ��E�����   �M��t��tVQP���  ���u؋���Q���  �htS��hP  V�Ѓ��E���tP��t��tVWP��  ���M����+���RH��PQ�E���   S�Ѓ���u�M�Q��  �U�R��  ��_^3�[��]á���HH���   j h�  S�҉E�����HH���   j h(  S��3�3���3��E��}ĉ]�9]��:  �U��څ��  �E�    ����   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T�Y�Z�Y �Z�Y$�Z�Y(�R�]��Q,�U�@����0��;�|��}ă|� �t   �U��M�ύI�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�Tv�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}�C�]�;]�������M�3�3�;�~�U���$    �t���   @;�|��U�R�  ���E�P��  ��_^�   [��]�˕ Օ �� � ������������U��E� �M+]� ���������������U��V��V�dS����Hl�AR�Ѓ��Et	V��  ����^]� ���������̋�� �S����������S���������̅�t��j�����̡���P��  �����P��(  ��U�����P��   ��V�E�P�ҋuP���zA  �M��A  ��^��]� ��������̡���P��$  ��U�����H��  ]��������������U�����H���  ]�������������̡���H��  ��U�����H���  ]��������������U�����H��x  ]��������������U�����H��|  ]��������������U���EV����St	V�H  ����^]� �������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V��迆  �����   �ESP�M��?  ����Q�J�E�P�ы���B�Pj j��M�h�SQ�҃��E�P�M���>  j j��M�Q�U�R��d���P�4Q  ��P�M�Q��B  ��P�U�R�B  ���P�߇  ���M����?  �M���>  ��d�����>  �M���>  ����H�A�U�R�Ѓ��M���>  ��[t	V��  ����^��]� ���U��EVP���q�  �����^]� �����Q躅  Y���������U��E�M�U�H4�M�P �U��M�@� �@8�y�@< � �@@�y�@D`y�@H�y�@L� �@Ppy�@l � �@X�y�@\Р �@`@� �@d� �@TP� �@h0� �@p�� �@t� �P0�H(�@,    ]��������������U���   h�   ��`���j P���  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj蕖����8��]��������������̋�`<����������̋�`0����������̋�`@����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`(����������̋�`8����������̋�`�����������U��V�u���t����QP��Ѓ��    ^]���������̡���H��@  hﾭ���Y����������U��E��t����QP��@  �Ѓ�]����������������U�����H���  ]��������������U�����H��  ]�������������̡���H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�r�  ������u_^]Ã} tWj V���  ��_������F��   ^]���U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW���  ������u_^]�Wj V�f�  ��_������F��   ^]�������������U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�v�  ������u_^]�Wj V���  ��_������F��   ^]�������������U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW���  ������u_^]�Wj V�f�  ��_������F��   ^]�������������U�����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�v�  ������u_^]�Wj V���  ��_������F��   ^]�������������U��M��t-�=� t�y���A�uP��  ��]á���P�Q�Ѓ�]��������U��M��t-�=� t�y���A�uP�l�  ��]á���P�Q�Ѓ�]��������U�����H�U�R�Ѓ�]���������U�����H�U�R�Ѓ�]���������U�����E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�2�  ������u_^]�Wj V��  ��_������F��   ^]���������U�����E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]Ã�s�   VW�xW��  ������u_^]Ã} tWj V���  ��_������F��   ^]����������U��E��u�   �����t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��  ������u_^]�Wj V�s�  ��_������F��   ^]����������U��E��u�   �����t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�p�  ������u_^]�Wj V���  ��_������F��   ^]�������U�����H�U�R�Ѓ�]���������U�����H�U�R�Ѓ�]���������U�����H�U�R�Ѓ�]���������U�����H�U�R�Ѓ�]���������U�����Hp�]�����Hp�h   �҃�������������U��V�u���t����QpP�B�Ѓ��    ^]���������U�����Pp�EP�EPQ�J�у�]� U�����Pp�EP�EPQ�J�у�]� U�����Pp�EP�EPQ�J�у�]� U�����Pp�EPQ�J�у�]� ���̡���HL���   ��U�����H@�AV�u�R�Ѓ��    ^]�������������̡���HL�������U�����H@�AV�u�R�Ѓ��    ^]�������������̡���PL���   Q�Ѓ�������������U�����PL�EP�EPQ���   �у�]� �������������U����V��HL���   V�҃���u����U�HL���   j RV�Ѓ�^]� ������   �ȋBP�Ћ�����   �MP�BH��^]� �����̡���PL��(  Q�Ѓ�������������U�����PL�EP�EPQ��,  �у�]� ������������̡���HL�Q�����U�����H@�AV�u�R�Ѓ��    ^]��������������U�����PL�E�R��VPQ�M�Q�ҋu��P���(  �M��(  ��^��]� ����U�����PL�EPQ���   �у�]� �U�����PL�EP�EPQ�J�у�]� ����PL�BQ�Ѓ���������������̡���PL�BQ�Ѓ���������������̡���PL�BQ�Ѓ����������������U�����PL�EP�EP�EPQ�J �у�]� ������������U�����PL�EPQ��4  �у�]� �U�����PL�EP�EP�EPQ�J$�у�]� ������������U�����PL�EP�EP�EP�EPQ�J(�у�]� �������̡���PL�B,Q�Ѓ���������������̡���PL�B0Q�Ѓ����������������U�����PL�EP�EPQ��  �у�]� ������������̡���PL���   Q�Ѓ�������������U�����PL�E��  ��VPQ�M�Q�ҋu��P���&  �M��&  ��^��]� ̡���PL�B4Q�Ѓ���������������̡���PL�B8j Q�Ѓ��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL���   ]��������������U�����PL�EPQ�J<�у�]� ���̡���PL�BQ��Y�U�����PL�EP�EPQ�J@�у�]� U�����PL�Ej PQ�JD�у�]� ��U�����PL�Ej PQ�JH�у�]� ��U�����PL�EjPQ�JD�у�]� ��U�����PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���T�  ���M����g�����t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �N���j�M�Q�U�R��轊  �M�赱��������   ��U�R�Ѓ�^��]�����������U���$����UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��ʾ��j�E�P�M�Q���9�  �M��1���������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��J���j�E�P�M�Q��蹉  �M�豰��������   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���4�  ���M����G�����t+�u���Y+  ������   ��U�R�Ѓ�_��^[��]� ������   �JL�E�P�ыu��P����+  ������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��$���W�M�Q�U�R���t�  ���M���臯����t+�u���*  ������   ��U�R�Ѓ�_��^[��]� ������   �JL�E�P�ыu��P���+  ������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��d���W�M�Q�U�R��贇  ���M����Ǯ��_^��[t������   ��U�R�������]Ë�����   �J<�E�P���]�������   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}�贻��W�M�Q�U�R����  ���M���������t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���T�  ���M����g�����t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� �����̡���PL���   Q��Y��������������U�����PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U�����PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��t���W�M�Q�U�R���Ą  ���M����׫����t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�褸��W�M�Q�U�R����  ���M���������t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��Է��W�M�Q�U�R���$�  ���M����7�����t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���T�  ���M����g�����t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �O���j�M�Q�UR��辁  �M趨��������   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��ߵ��j�U�R�E�P���N�  �M��F���������   �
�E�P�у�^��]� ��������U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��Z���j�E�P�M�Q���ɀ  �M������������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��ڴ��j�E�P�M�Q���I�  �M��A���������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��Z���j�E�P�M�Q����  �M������������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��ڳ��j�E�P�M�Q���I  �M��A���������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��o���j�U�R�E�P����~  �M��֥��������   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���T~  ���M����g�����t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��4���W�M�Q�U�R���}  ���M���藤����t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}�脱��W�M�Q�U�R����|  ���M���������t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}�蚰��j�E�P�M�Q���	|  �M�����������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��/���j�U�R�E�P���{  �M�薢��������   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�迯��j�U�R�E�P���.{  �M��&���������   �
�E�P�у�^��]� ��������U�����H���   ]��������������U�����H���   ]�������������̡���H���   �����H���   ��U�����H���   V�u�R�Ѓ��    ^]�����������U�����H���   ]��������������U�����HL�QV�ҋ���u^]á���H�U�ER�UP���  RV�Ѓ���u����Q@�BV�Ѓ�3���^]����������U�����H�U�E���  R�U�� P�ERP�у�]������U�����H���   ]��������������U�����H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡���PL�BLQ�Ѓ���������������̡���PL�BPQ�Ѓ����������������U�����PL�EP�EPQ�JT�у�]� U�����PL�EPQ��  �у�]� �U�����PL�EPQ���   �у�]� ̡���PL�BXQ�Ѓ����������������U�����PL�EP�EP�EPQ�J\�у�]� ������������U���4���SV��HL�QW�ҋ�3ۉ}�;��x  �M��  ����E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�����   �BSSW���Ѕ���   ����QL�BW�Ћ���;���   ��    ������   �B(���ЍM�Qh�   ���u��u��������   �M�;���   ������   ���   S��;�tm������   �ȋB<V�Ћ�����   ���   �E�P�у�;�t����B@�HV�у���;��\����}��M������M���  ��_^[��]� �}�����B@�HW�ы�����   ���   �M�Q�҃��M��Ɋ���M��  _^3�[��]� �����̡���PL�B`Q�Ѓ���������������̡���PL�BdQ�Ѓ����������������U�����PL�EPQ�Jh�у�]� ���̡���PL��D  Q�Ѓ������������̡���PL�BlQ�Ѓ����������������U�����PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh`� h@� h � h� R�Q�U R�UR�UR�U���A�$�5���vLRP���   Q�Ѓ�4^]�  ������̡���PL���   Q�Ѓ�������������U�����PL�EP�EP�EPQ��   �у�]� ���������U�����PL��H  ]�������������̡���PL��L  ��U�����PL��P  ]��������������U�����PL��T  ]��������������U�����PL�EP�EP�EP�EP�EPQ���   �у�]� �U�����PL�EP�EP�EPQ���   �у�]� ���������U�����PL�EP�EP�EP�EPQ��   �у�]� �����U�����HL���   ]��������������U�����HL���   ]��������������U�����HL���   ]�������������̡���HL��  �����HL��@  ��h�Ph^� ��5  ���������������U��Vh�j\h^� ���5  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� ���V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\����QLjP���   ���ЋM��U�Rh=���M�}��p����������   ���   �U�R�Ѓ��M��u��\�����_^��]Ë�����   ���   �E�P�у��M��u��.���_�   ^��]����U��� ���V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\����QLjP���   ���ЋM��U�Rh<���M�}���o����������   ���   �U�R�Ѓ��M��u�茅����_^��]Ë�����   ���   �E�P�у��M��u��^���_�   ^��]���̡��V�񋈈   ���   V�҃��    ^���������������� �������������U���d�}W��t�   _��]� ���Pt�U�S�U�]�]�S�҉E��u[�   _��]� ����U�HH��   VRS�Ћ���Qd�J<�E��EP�эU�j/R���Bp���E�jP�7p������Qd�E�JpVSP�у�(3�j ��u����Bd�U�@�M�QR�������Qd�M�R�E�PQ��3���9u~a3�;u���;�uO�E��RxVP�M�Q����� �U��@�]��@�]���S����t����Hd�E���   j j�U�RP�у�F;u|�C���W���^[�   _��]� �������U����E�P�P�]� �������������  �������������3�� �����������U����   �ES��t
���[��]� ����PH�M�R,VW��$���P�ҋ���Pt�   �}��}W���E�����3��҅���   ���PxVW�M�Q����� �@�@��S������A�|   �E�����ˋUR�U��E����M����E������]��E����E��E������E������]��E������E��E������E������]�Hd�E�IP�ERP�у���t�E�u�t������؋�BtW��F��;��A����E�_^[��]� �����U������SVW�}��H@�Q8j W�ҋ]��Rx��SW�M�Q���ҋE�@��E�R|�Ƀ��ɋ�� �@0�E��������@H�E��������@ ���@�@8�����@P�����@(�����@�@@�����@X����S����������X�X�EP��_^�   [��]� ���������3�� �����������3�� ����������̸   �$ ��������� �������������� �������������� �������������3�� �����������3�� �����������U��UP�EQWRPV���������   ǆ�   �yǆ�   �yǆ�   Pyǆ�   `� ǆ�   �� ǆ�   �� ǆ�   @� ]������������U�����P�B<��   V�u���Ѕ�t�Mj VQ�T�������u^��]�SWh   ������j R裹  �]�E�}�M SP3��������(������E��� ��t�E��� �� t�E��� ��y�E�P� _��[t�E�p� �U�Eh   ������QRPj�h����^��]����������̋�`\����������̋�`l����������̋�`P����������̋�``����������̋�`p����������̋�`T����������̋�`d����������̋�`X����������̋�`h����������̡���H\�������U�����H\�AV�u�R�Ѓ��    ^]�������������̡���P\�BQ�Ѓ���������������̡���P\�BQ�Ѓ����������������U�����P\�EPQ�J�у�]� ����U�����P\�EP�EPQ�J�у�]� U�����P\�EPQ�J�у�]� ���̡���P\�BQ�Ѓ����������������U�����P\�EPQ�J �у�]� ����U�����P\�EP�EPQ�J$�у�]� U�����P\�EP�EP�EPQ�J(�у�]� ������������U�����P\�EPQ�J0�у�]� ����U�����P\�EPQ�J@�у�]� ����U�����P\�EPQ�JD�у�]� ����U�����P\�EPQ�JH�у�]� ���̡���P\�B4Q�Ѓ����������������U�����P\�EP�EPQ�J8�у�]� U�����P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu���#  ����H\�QV�҃���S����#  3���~=��I ����H\�U�R�U��EP�A(VR�ЋM��Q���#  �U�R���#  F;�|�_^[��]� ���������������U���VW�}�E��P����  �}� ��   ����Q\�BV�Ѓ��M�Q����  �E���t]S3ۅ�~H�I �UR���  �E�P���  �E;E�!������Q\P�BV�ЋE@���E;E�~�C;]�|�[_�   ^��]� _�   ^��]� ����P�BVj j����Ћ�^���������U�����P�E�RVj P���ҋ�^]� U�����P�E�RVPj����ҋ�^]� ����P�B�����U�����P���   Vj ��Mj V�Ћ�^]� �����������U�����P�EPQ�J�у�]� ����U�����P�EPQ�J�у����@]� ���������������U�����P�E�RtP�ҋ�����   P�BX�Ѓ�]� ���U�����P�E�Rlh#  P�EP��]� ���������������U�����P�E�RlhF  P�EP��]� ���������������U�����P�E�RtP�ҋ�����   �M�R`QP�҃�]� ���������������U�����P���   ]��������������U�����P�E���   P�҅�u]� ������   P�B�Ѓ�]� �������̡���PD�BQ�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�BQ�Ѓ����������������U�����PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U�����PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�����PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�����PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U�����PX�EPQ�J�у�]� ����U�����PX�EPQ�J�у�]� ����U�����PX�EPQ�J�у�]� ����U�����PX�EPQ�J�у�]� ����U�����PX�EPQ�J$�у�]� ����U�����PX�EPQ�J �у�]� ����U�����PD�EP�EPQ�J�у�]� U�����HD�U�j R�Ѓ�]�������U�����H@�AV�u�R�Ѓ��    ^]��������������U�����HD�	]��U�����H@�AV�u�R�Ѓ��    ^]��������������U�����HD�U�j R�Ѓ�]�������U�����H@�AV�u�R�Ѓ��    ^]��������������U�����U�HD�Rh'  �Ѓ�]����U�����H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h�  �҃�����������U�����H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h:  �҃�����������U�����H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E�������   �R�E�Pj�����#E���]�̡���HD�j h�F �҃�����������U�����H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h�_ �҃�����������U�����H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E�����E�    ���   �R�E�Pj������؋�]� ̡���PD�B$Q�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡��V��H�QV�ҡ���H$�QDV�҃���^�����������U����V��H�QV�ҡ���H$�QDV�ҡ���U�H$�AdRV�Ѓ���^]� ��U����V��H�QV�ҡ���H$�QDV�ҡ���U�H$�ARV�Ѓ���^]� ��U����V��H�QV�ҡ���H$�QDV�ҡ���H$�U�ALVR�Ѓ���^]� �̡��V��H$�QHV�ҡ���H�QV�҃�^�������������U�����P$�EPQ�JL�у�]� ����U�����P$�R]�����������������U�����P$�Rl]����������������̡���P$�Bp����̡���P$�BQ�Ѓ����������������U�����P$��VWQ�J�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]� ���U�����P$�EPQ�J�у�]� ����U�����P$��VWQ�J �E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]� ���U�����P$��VWQ�J$�E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]� ���U���,VW�E�P�o�������Q$�JP�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у� _��^��]� �����̡���P$�B(Q��Yá���P$�BhQ��Y�U�����P$�EPQ�J,�у�]� ����U�����P$�EPQ�J0�у�]� ����U�����P$�EPQ�J4�у�]� ����U�����P$�EPQ�J8�у�]� ����U�����UV��H$�ALVR�Ѓ���^]� ��������������U�����H�QV�uV�ҡ���H$�QDV�ҡ���H$�U�ALVR�Ћ���E�Q$�J@PV�у���^]�U�����UV��H$�A@RV�Ѓ���^]� ��������������U�����P$�EPQ�J<�у�]� ����U�����P$�EPQ�J<�у����@]� ���������������U�����P$�EP�EPQ�JP�у�]� U�����P$�EPQ�JT�у�]� ���̡���H$�QX�����U�����H$�A\]�����������������U�����P$�EP�EP�EPQ�J`�у�]� �����������̡���H(�������U�����H(�AV�u�R�Ѓ��    ^]��������������U�����P(�R]����������������̡���P(�B�����U�����P(�R]�����������������U�����P(�R]�����������������U�����P(�R ]�����������������U�����P(�E�RjP�EP��]� ��U�����P(�E�R$P�EP�EP��]� ����P(�B(����̡���P(�B,����̡���P(�B0�����U�����P(�R4]�����������������U�����P(�RX]�����������������U�����P(�R\]�����������������U�����P(�R`]�����������������U�����P(�Rd]�����������������U�����P(�Rh]�����������������U�����P(�Rx]�����������������U�����P(�Rl]�����������������U�����P(�Rt]�����������������U�����P(�Rp]�����������������U�������E�    �E�    �P(�RhV�E�P���҅���   �E���uG����H�A�U�R�Ћ���Q�E�RP�M�Q�ҡ���H�A�U�R�Ѓ��   ^��]� ����Qh�Sh8  P���   �Ћ�����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�ֺ����3�^��]� ����E��Q�M�j HP�EQ�JP�эU�R褺�����   ^��]� �����U������V��H�A�U�R�Ѓ��M�Q������^��u����B�P�M�Q�҃�3���]� ����H$�E�I�U�RP�ы���B�P�M�Q�҃��   ��]� �U��Q����P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U�����P(�R8]�����������������U�����P(�R<]�����������������U�����P(�R@]�����������������U�����P(�RD]�����������������U�����P(�RH]�����������������U�����P(�E�R|P�EP��]� ����U�����P(�RL]�����������������U�����E�P(�BT���$��]� ���U�����E�P(�BPQ�$��]� ����̡���H(�Q�����U�����H(�AV�u�R�Ѓ��    ^]��������������U�����P(���   ]��������������U�����H(�A]����������������̡���H,�Q,����̡���P,�B4�����U�����H,�A0V�u�R�Ѓ��    ^]�������������̡���P,�B8�����U�����P,�R<��VW�E�P�ҋu������H�QV�ҡ���H$�QDV�ҡ���H$�QLVW�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у�_��^��]� �������U�����P,�E�R@��VWP�E�P�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ��̡���H,�j j �҃��������������U�����P,�EP�EPQ�J�у�]� U�����H,�AV�u�R�Ѓ��    ^]�������������̡���P,�B����̡���P,�B����̡���P,�B����̡���P,�B ����̡���P,�B$����̡���P,�B(�����U�����P,�R]�����������������U�����P,�R��VW�E�P�ҋu������H�QV�ҡ���H$�QDV�ҡ���H$�QLVW�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у�_��^��]� �������U�����H��D  ]��������������U�����H��H  ]��������������U�����H��L  ]��������������U�����H�I]�����������������U�����H�A]�����������������U�����H�I]�����������������U�����H�A]�����������������U�����H�I]�����������������U�����H���  ]��������������U�����H�A]�����������������U���V�u�E�P���+�������Q$�J�E�P�у���u-����B$�PH�M�Q�ҡ���H�A�U�R�Ѓ�3�^��]Ë���Q�J�E�jP�у���u=�U�R��������u-����H$�AH�U�R�Ћ���Q�J�E�P�у�3�^��]Ë���B�HjV�у���u����B�HV�у����I�������Q$�JH�E�P�ы���B�P�M�Q�҃��   ^��]�����������U�����H�A ]�����������������U�����H�I(]�����������������U�����H��  ]��������������U�����H��   ]��������������U�����H��  ]��������������U�����H��  ]��������������U�����H�A$��V�U�WR�Ћ���Q�u���BV�Ћ���Q$�BDV�Ћ���Q$�BLVW�Ћ���Q$�JH�E�P�ы���B�P�M�Q�҃�_��^��]������U�����H���  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q$�BDV�Ћ���Q$�BLVW�Ћ���Q$�JH�E�P�ы���B�P�M�Q�҃�_��^��]���U�����H���  ]��������������U���<���SVW�E�    ��t�E�P�   �������/����Q�J�E�P�   �ы���B$�PD�M�Q�҃��}����H�u�QV�ҡ���H$�QDV�ҡ���H$�QLVW�҃���t)����H$�AH�U�R����Ћ���Q�J�E�P�у���t&����B$�PH�M�Q�ҡ���H�A�U�R�Ѓ�_��^[��]���U�����H�U���  ��VWR�E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡���H���   ��U�����H���   V�uV�҃��    ^]�������������U�����P�]�����P�B����̡���P���   ��U�����P�R`]�����������������U�����P�Rd]�����������������U�����P�Rh]�����������������U�����P�Rl]�����������������U�����P�Rp]�����������������U�����P�Rt]�����������������U�����P���   ]��������������U�����P�Rx]�����������������U�����P���   ]��������������U�����P�R|]�����������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P�EPQ��  �у�]� �U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U��E��t ����R P�B$Q�Ѓ���t	�   ]� 3�]� U�����P �E�RLQ�MPQ�҃�]� U��E��u]� ����R P�B(Q�Ѓ��   ]� ������U�����P�R]�����������������U�����P�R]�����������������U�����P�R]�����������������U�����P�R]�����������������U�����P�R]�����������������U�����P�R]�����������������U�����P�E�R\P�EP��]� ����U�����E�P�B ���$��]� ���U�����E�P�B$Q�$��]� �����U�����E�P�B(���$��]� ���U�����P�R,]�����������������U�����P�R0]�����������������U�����P�R4]�����������������U�����P�R8]�����������������U�����P�R<]�����������������U�����P�R@]�����������������U�����P�RD]�����������������U�����P�RH]�����������������U�����P�RL]�����������������U�����P�RP]�����������������U�����P���   ]��������������U�����P�RT]�����������������U�����P�EPQ��  �у�]� �U�����P���   ]��������������U�����P���   ]��������������U�����P�RX]����������������̡���P���   ��U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]��������������U�����P���   ]�������������̡���P���   ��U�����P���   ]�������������̡���P���   �����P���   �����P���   ��U�����H���   ]��������������U�����H��   ]��������������U�����H�U�E��VWRP���  �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]������������U�����H���  ]��������������U�����P(�} �R8����P��]� �U�����P�BdS�]VW��j ���Ћ���Qh�S�p���   hc  V�Ћ�����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ���Q(�BHV���Ѕ�t ����Q(�E�R VP���҅�t�   �3��EP������_��^[]� ������U�����U�� V��H$�IWR�E�P�ы�����B�P�M�Q�ҡ���H�A�U�RW�Ћ���Q�J�E�P�у��U�R������������H�A�U�R�Ѓ�_��^��]� �����������U�������   �BXQ�Ѓ���u]� ����Q|�M�RQ�MQP�҃�]� ���U�������   �BXQ�Ѓ���u]� ����Q|�M�R8Q�MQP�҃�]� ���U��EV��j �����Qj j P�B�ЉF����^]� ��̡��Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ����Q�MP�EP�Q�JP�у��F�   ^]� ����U��E�M�UP��P�EjP�>����]��������������̸   �����������U��V�u��t���u6�EjP�>������u3�^]Ë��?����t���t��U3�;P��I#�^]�������U��� �E�M���  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��4�E��}���t�u+��\�P@�M���u�EH�E����   )}��u��	;]��u��s���u�]�;]}�M��>P�E�V�Ѕ�y�u�C�]�M��E��VP�҅��d����F��}��t�M�+���I ��P@�M��T�u�]��;]~��/���_^[��]� ������U���(W�}�����E�E�M���/  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��
�U���$    ��~�M�M�J)}��U��G�M�E��M��t'�M�+����$    ��pf�\���M�f�f�4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��H����}�F���t!�M�+ȍI �Pf���Of�f�T�u�]��}�;E�~����	���^[_��]� ����������U���(W�}�����E�E�M���  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��9�M�E��M��t�M�+ȋ\�p���M��4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��W����}�F���t�M�+Ȑ��P��O��T�u�]��}�;E~��"���^[_��]� ��U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   xO�E�   �}��}_^3�[��]� �}}���E������uu��VP�҅�tyO�}�G�}��E9E�~�_^3�[��]� ��~3�E���]��]�E����E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   y�M_^�    3�[��]� �O�3��E�   �M��} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�ty�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �����������������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH������������Dz�u�؋��3�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�����U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� ��3ɉ�H�H�H�V��V�'����FP����3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}��'	  S�]����  ��؋���M�U��>���U�@�U���� �U��@�@�B�@�������@���@�   ���]��E��U�;���  �w�����  �w�������F�܍B��   �U������������ˋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]����]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]��]��U���E��U��R�э����N�B���B�P���R���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]�����B���B���U����E��������]��E����E����������E������E��E��U����E��]����E��U��E��U��T����E�ɋU�����������;���   �ߍ���+�������͋�@�������O�]��@���]��@���U������M������]��E��E����E������E����������E��E��U����E��]����E��U��E��E��U�u�������������������������[�[�E����������������s  ��������������Dz���������E��+������������������M����M��E������������������[H���[P���[X�E����E���������zu������������zh�����CP���CX���CH���CX�������cH���[���[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@��   ������������z]�CX���CP�����cH�CH���CP�������[�[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@�]�CP���CX�����CH���CX�����cP���[0���[8�[@�C8�KX�C@�KP���CH�K@�C0�KX���C0�KP�C8�KH�����[�[ �[(��$���SQ�����E��U�   �����}��M������3�3��u��u���|)�A�����B�4�u�0u��u�p��J�u�u�U�E;�}�Q���E���u��U��1���@���K�I�E    ��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]�� �K��C0�H���@�KH��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���U����n  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������]��E�E����]���E����]��E��M����@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������U��E��]��E��U������������������9M|��[��_��^���؋�]� ���������ʋE�����׋��@�E�Ѝ��K��C0�H���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���CX�H�E@�E���]����E��������������������M����������]��E��E�;��T�����[������_��^��]� �����h�Ph_� �������������������h�jh_� �o�������uË@����U��V�u�> t/h�jh_� �C�������t��U�M�@R�Ѓ��    ^]���U��Vh�jh_� ���	�������t�@��t�MQ����^]� 3�^]� �������U��Vh�jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh�jh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�jh_� ���9�������t�@��t�MQ����^]� 3�^]� �������U��Vh�j h_� �����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�j$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh�j(h_� ���|�������t�@(��t��^��3�^������Vh�j,h_� ���L�������t�@,��t��^��3�^������U��Vh�j0h_� ����������t�@0��t�MQ����^]� 3�^]� �������U��Vh�j4h_� �����������t�@4��t�M�UQR����^]� ���^]� ��Vh�j8h_� ����������t�@8��t��^��3�^������U��Vh�j<h_� ���i�������t�@<��t�MQ����^]� ��������������U��Vh�j@h_� ���)�������t�@@��t�MQ����^]� ��������������U��Vh�jDh_� �����������t�@D��t�MQ����^]� 3�^]� �������U��Vh�jHh_� ����������t�@H��t�MQ����^]� ��������������Vh�jLh_� ���l�������t�@L��t��^��3�^������Vh�jPh_� ���<�������t�@P��t��^��3�^������Vh�jTh_� ����������t�@T��t��^��^��������Vh�jXh_� �����������t�@X��t��^��^��������Vh�j\h_� ����������t�@\��t��^��^��������U��Vh�j`h_� ���y�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�jdh_� ���9�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh�jhh_� �����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�jlh_� ����������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�jph_� ���Y�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�jth_� ����������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�jxh_� �����������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh�j|h_� ����������t�@|��t�MQ����^]� 3�^]� �������U��Vh�h�   h_� ���V�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�h�   h_� ���F�������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������M�������_�U�^��[�U����U��������������������c  ��������������D�Ez���P�P���]� �������E�����E����X�M��X��]� ����U���@��S�A���E�    �����]����]��]�� T�������]����]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P������F�@��R�M������~���Q�M������v;�t�v��P�M������M����M��M�u��}� _^[tV�E؋E�E����E��E����E��E����T������������X���X��� ���`���`�E����X�X��]� ��E����������P���P�E����X�X��]� �����������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��x+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~!V�1�d$ ���   @u	�����t@��Ju�^�����̋QV3���~�	�d$ ����ШtF��Ju��^�����������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%����E���;�}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$���E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��2H[o�����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP����3����F�F^��U��SV��WV�����^S�����E3����~�~;�t_����Q���   hT��jIP�у��;�t9�}��t;����B���   hT��    jNQ�҃����uV�{�����_^3�[]� �E�~_�F^�   []� ����������U��V��WV�C����FP�:����}���F    �F    ����   �? ��   �G����   ����Q���  hT��jlP�у����t>� t@�G��t9����JhT��    ���  jqR�Ѓ��F��u���v���_3�^]� �O��N�G�F��    ���t��t��tQPR�d  ���F��t�VP��RP�GP�  ��_�   ^]� ��������U��SV��WV�2����~W�)���3����F�F9E�  �];���   ����QhT��    h�   P���  �Ѓ����t@�} tN�]��tD����Q���  hT��    h�   P�у����u���n���_^3�[]� �^�]�0�]�F   ����B���  hTh�   j�у����t���^��t��    ��t�UQRP��b  ���E��t!�N�?�W�QWP�R  ��_^�   []� ��_^�   []� ���U��Q�A�E� ��~JS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U���Ou�_^[�E��Ћ�]� �����������U��S�]V��3�W�~���F�F�CV;C��   �d~��W�^~��3��F�F����Q���   hTjIj�Ѓ������   ����Q���   hTjNj�Ѓ����uV�~����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� ��}��W�}��3��F�F����B���   hTjIj�у����t[����B���   hTjNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�@`  ��]�����������̡���H���   ��U�����H���   V�u�R�Ѓ��    ^]����������̡���P���   Q�Ѓ�������������U�����P�EPQ���   �у�]� ̡���H�������U�����H�AV�u�R�Ѓ��    ^]��������������U�����H�AV�u�R�Ѓ��    ^]��������������U�����P��Vh�  Q���   �E�P�ы�����   �Q8P�ҋ������   ��U�R�Ѓ���^��]��������������̡���P�BQ�Ѓ����������������U�����P�EPQ�J\�у�]� ����U�����P�EP�EP�EP�EP�EPQ���   �у�]� �U�����P�EP�EP�EP�EPQ�JX�у�]� �������̡���P�B Q��Y�U�����P�EP�EP�EP�EPQ���   �у�]� �����U�����P�EP�EP�EPQ�J�у�]� ������������U�����H��   ]��������������U�����P�R$]�����������������U�����P�EP�EP�EP�EPQ�J(�у�]� ��������U�����P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U�����P�EP�EP�EP�EPQ�J,�у�]� ��������U����V��H�QWV�ҍx�����H�QV�ҋ���Q�M�R4Q�MQ�MQWHPj j V�҃�(_^]� ���������������U�����P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U�����P�EP�EPQ�J@�у�]� U�����P�EPQ�JD�у�]� ���̡���P�BLQ�Ѓ���������������̡���P�BLQ�Ѓ���������������̡���P�BPQ�Ѓ����������������U�����P�EPQ�JT�у�]� ����U�����P�EPQ�JT�у�]� ����U�����P�EP�EPQ���   �у�]� �������������U�����P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у� ��^��]� ������̡���P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡���H�������U�����H�AV�u�R�Ѓ��    ^]��������������U�����P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�����P�EPQ�J�у�]� ���̡���P�BQ��Y�U�����P�EP�EPQ�J�у�]� U��VW���p���M�U�x@�EPQR���p���H ���_^]� �U��VW���tp���M�U�xD�EPQR���^p���H ���_^]� �V���Hp���xH u3�^�W���6p���΍xH�,p���H �_^�����U��V���p���xL u3�^]� W��� p���M�U�xL�EPQR����o���H ���_^]� �������������U��V����o���xP u���^]� W���o���M�U�xP�EP�EQRP���o���H ���_^]� ��������U��V���uo���xT u���^]� W���_o���M�xT�EPQ���Mo���H ���_^]� U���S�]VW���t.�M��f������o���xL�E�P���o���H ��ҍM�蠦���}��tZ����H�A�U�R�Ћ���Q�J�E�WP�ы���B�P�M�Q�҃����n���@@��t����QWP�B�Ѓ�_^[��]� ������U��VW���n���xH�EP���vn���H ���_^]� ���������U��VW���Tn���M�U�xD�EP�EQRP���:n���H ���_^]� �������������U��V���n���xP u
�����^]� W����m���M�U�xP�EP�EQ�MR�UPQR����m���H ���_^]� ��������������U��V���m���xT u
�����^]� W���m���M�xT�EPQ���m���H ���_^]� ��������������U��V���em���xX tW���Wm���xX�EP���Im���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��(5  ����t.�E�;�t'����J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡���H��   ��U�����H��$  V�u�R�Ѓ��    ^]�����������U�����UV��H��(  VR�Ѓ���^]� �����������U�����P�EQ��,  P�у�]� �U�����P�EQ��,  P�у����@]� �����������̡���H��0  �����H��4  ��U��E��t�@�3�����RP��8  Q�Ѓ�]� �����U�����P�EPQ��<  �у�]� �U�����P�EP�EP�EPQ��@  �у�]� ���������U�����P�EP�EPQ��D  �у�]� �������������U�����P�EPQ��H  �у�]� �U�����P�E��L  ��VWPQ�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ��������������̡���P��T  Q�Ѓ������������̡���P��P  Q�Ѓ�������������U�����P�EPQ��X  �у�]� ̡���H��\  ��U�����H��`  V�u�R�Ѓ��    ^]�����������U�����P�EP�EP�EP�EP�EPQ��d  �у�]� �U�����P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���O褪����3��G �G$�G(�G,�G0�G4�G8�G<�G@�GD�GH�GL�GP�GT�GX�G\�_p��G`�Gd�Gh�Gx�����G|   ��_^����������������V��W�>��t7���i���xP t$S���i��j j �XPj�FP����h���H ���[�    �~` t����H�V`�AR�Ѓ��F`    _^������������U��SV��Fx����Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�������u#���hPT����H��0  h�   �҃��E�~P��蜭���j j jW�N����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ����Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��QV��~d tg�E;Fxt_�N`W�>�M����kg���xP u����(S���Xg���UR�XP�E�Pj�NQ���@g���H ���[�F|_��u�E�Fx�E��t�    �F`^��]� �M�Fx������t�3�^��]� ���������U��QVW�}����1  ����H�QhV�҃������u"�H��0  hPTh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���?/  �EF;u�|�UR�k����_�   ^��]� �������������U��QVW�}�����0  ����H�QhV�҃������u"�H��0  hPTh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'������QP�Bh�Ѓ���t�M��R���\.  F;u�|ʍEP�j����_�   ^��]� �������������hPTh�   h�h�   �wn������t������3��������V��������N^�������������������U��VW�}�7��t�������N����V�]m�����    _^]Ë�3ɉH��H�@   �������������U��ыM��tK�E��t������   P�B@��]� �E��t������   P�BD��]� ������   R�PD��]� �����U�����P@�Rd]�����������������U�����P@�Rh]�����������������U�����P@�Rl]�����������������U�����P@�Rp]�����������������U�������   ���   ]�����������U�������   ���   ]����������̡���P@�Bt����̡���P@�Bx�����U�����P@�R|]����������������̡���P@���   �������   �Bt��U�����P@���   ]�������������̡���P@���   ��U�����P@���   ]��������������U�����P@���   ]��������������U�����P@���   ]��������������U�����P@���   ]��������������U����V��H@�QV�ҋM����t��#�������Q@P�BV�Ѓ�^]� �̡���PH���   Q�Ѓ�������������U�����P@�EPQ�JL�у�]� ���̡���P@�BHQ�Ѓ����������������U�����P@�EP�EP�EPQ�J�у�]� ������������U�����P@�EPQ�J�у�]� ����U�����P@�EP�EPQ�J�у�]� U�����P@�EPQ�J �у�]� ����U�������   �R]��������������U�������   �R]��������������U�������   �R ]��������������U�������   ���   ]�����������U�������   ��D  ]�����������U�����E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U�������   ���   ]����������̡�����   �B$�����H@�Q0�����U�����H@�A4j�URj �Ѓ�]����U�����H@�A4j�URh   @�Ѓ�]�U�����H@�U�E�I4RPj �у�]�̡���H|�������U��V�u���t����Q|P�B�Ѓ��    ^]��������̡���H|�Q �����U��V�u���t����Q|P�B(�Ѓ��    ^]��������̡���H@�Q0�����U��V�u���t����Q@P�B�Ѓ��    ^]���������U�����H@���   ]��������������U��V�u���t����Q@P�B�Ѓ��    ^]��������̡���PH���   Q�Ѓ�������������U�����PH�EPQ��d  �у�]� �U�����H �IH]�����������������U��}qF uHV�u��t?������   �BDW�}W���Ћ���Q@�B,W�Ћ���Q�M�Rp��VQ����_^]����������̡���P@�BT�����U�����P@�RX]�����������������U�����P@�R\]����������������̡���P@�B`�����U�����H��T  ]��������������U�����H@�U�A,SVWR�Ћ���Q@�J,���EP�ы���Z��h��hE  �΋������Ph��hE  ������P��T  �Ѓ�_^[]����h�Ph^� �`������������������U��Vh�jh^� ���9�������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh�jh^� �����������t�@��tV�Ѓ�^�3�^���U��Vh�jh^� ���ɽ������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh�jh^� ��能������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u��������N`��������   �������   ������ݞ�  ��^��]� ����U��Vh�jh^� �����������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh�jh^� ��蹼������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh�j h^� ���y�������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�j$h^� ���)�������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�j(h^� ����������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh�j,h^� ��註������t �@,�E���t�E�MPQV�U���^��]� ��^��]� ��������U��Vh�j0h^� ���Y�������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh�j4h^� ����������t�@4��tV�Ѓ�^�3�^���Vh�j8h^� ���ܺ������t�@8��tV�Ѓ�^�������U���`Vh�jDh^� ��覺������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u���������^��]� ����U��Vh�jHh^� ���I�������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh�jLh^� ���	�������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh�jPh^� ���ɹ������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh�jTh^� ��艹������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh�jXh^� ���I�������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh�j`h^� ����������t�@`��tV�Ѓ�^�3�^���U��Vh�jdh^� ��蹸������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh�jhh^� ���v�������t1�@h��t*�MQ�U�VR�Ћu��P����)���M�������^��]� �u�������^��]� �����������Vh�jph^� ����������t�@p��tV�Ѓ�^Ã��^��Vh�jlh^� ���ܷ������t�@l��tV�Ѓ�^Ã��^��Vh�jth^� ��謷������t�@t��tV�Ѓ�^�3�^���U��Vh�jxh^� ���y�������t�@x��t
�MQV�Ѓ�^]� ������������Vh�j|h^� ���<�������t�@|��tV�Ѓ�^�������Vh�h�   h^� ���	�������t���   ��tV�Ѓ�^�U��Vh�h�   h^� ���ֶ������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh�h�   h^� ��膶������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh�h�   h^� ���3�������tU���   ��tKW�M�VQ�Ћ���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]� ����H�u�QV�҃���^��]� ����������Vh�h�   h^� ��虵������t���   ��tV�Ѓ�^Ã��^������������U��Vh�h�   h^� ���V�������t���   ��t
�MQV�Ѓ�^]� ������U��Vh�h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h�   h^� ���ƴ������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh�h�   h^� ���y�������t���   ��tV�Ѓ�^�3�^�������������U��Vh�h�   h^� ���6�������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh�h�   h^� ��薳������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�h�   h^� ���F�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h�   h^� ��覲������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh�h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������Vh�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh�h�   h^� ���ٱ������t���   ��tV�Ѓ�^�3�^�������������Vh�h�   h^� ��虱������t���   ��tV�Ѓ�^�3�^�������������U��Vh�h�   h^� ���V�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh�h�   h^� ���	�������t���   ��tV�Ѓ�^�3�^�������������U���Vh�h�   h^� ���ð������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�h�   h^� ���F�������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�h�   h^� ���	�������t���   ��tV�Ѓ�^�3�^�������������U���Vh�h�   h^� ���ï������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�h�   h^� ���F�������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�h�   h^� ���	�������t���   ��tV�Ѓ�^�3�^�������������U��Vh�h�   h^� ���Ʈ������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh�h�   h^� ���u�������t#���   �E���t�E�MPQV�U���^��]� ��^��]� ��U��Vh�h�   h^� ���&�������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh�h�   h^� ���֭������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�h�   h^� ��膭������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h   h^� ���6�������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh�h  h^� ����������t��  ��tV�Ѓ�^�3�^�������������U���Vh�h  h^� ��裬������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�h  h^� ���#�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�h  h^� ��裫������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh�h  h^� ���&�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�h  h^� ����������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�h  h^� ��親������t��  ��t
�MQV�Ѓ�^]� ������Vh�h   h^� ���i�������t��   ��tV�Ѓ�^�3�^�������������U��Vh�h$  h^� ���&�������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h(  h^� ���֩������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h,  h^� ��膩������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�h0  h^� ���9�������t��0  ��tV�Ѓ�^�3�^�������������U��Vh�h4  h^� �����������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h8  h^� ��覨������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�h<  h^� ���V�������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh�h@  h^� ����������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�hD  h^� ��蹧������t��D  ��tV�Ѓ�^�3�^�������������U��Vh�hH  h^� ���v�������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�hL  h^� ���&�������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�hP  h^� ���֦������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh�hT  h^� ��腦������t'��T  �E���t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh�hX  h^� ���&�������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh�j<h^� ���٥������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh�j@h^� ��虥������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h�Ph�� �`������������������h�jh�� �?�������uË@����U��V�u�> t/h�jh�� ��������t��U�M�@R�Ѓ��    ^]���U��Vh�jh�� ���٤������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�jh�� ��艤������t�@��t�M�UQR����^]� ����������U��Vh�jh�� ���I�������t�@��t�M�UQR����^]� ����������U��Vh�jh�� ���	�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�j h�� ��蹣������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�j$h�� ���i�������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�j(h�� ����������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�j,h�� ���ɢ������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh�j0h�� ���i�������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�j4h�� ����������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh�j8h�� ��踡������t�@8�E���t�E�MPQ���U�^��]� ��^��]� ����������U��Vh�j<h�� ���i�������t�@<��t�M�UQR����^]� ����������U��Vh�j@h�� ���)�������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh�jHh�� ����������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh�jDh�� ��詠������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh�jLh�� ���h�������t#�@L�E���t�E�EP�����$�U�^��]� ��^��]� �����U��Vh�jPh�� ����������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh�jTh�� ���ٟ������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�jXh�� ��艟������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�j\h�� ���9�������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h�jh�� ��������t�@�ЉF�~��t6h�jh�� 軞������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h�jh�� �a�������t�@��t�M�UQR���Ѓ~ t1h�jh�� �0�������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h�jh�� ��������t�@�ЉF�v��t+h�jh�� 輝������t�@��t�M�UQR����^]� �������������U��V�q��t@h�jh�� �t�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h�j h�� ��������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h�jh�� ���������t�@�ЉF�}�]�M�UWSQR���  ��t;�v��t4h�j$h�� ��������t�@$��t�M�UWSQR����_^[]� _^3�[]� ���U��V�q��t8h�j(h�� �4�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��V�q��tHh�j,h�� ��������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  ������U��V�q��t<h�j0h�� 脛������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��EHu�E�M�������   ]� �������������U��EHV����   �$�dc�   ^]á �@� ���uT�EP�������=�.  }�����^]Ëu��t�h�Tjmh�j�B������t ���]z�������tV���~���   ^]����    �   ^]ËM�UQR�����������H^]�^]�0���� �u.�ӭ���^��������t����z��V�WA�������    �   ^]Ã��^]Àbc cxb^c�b����h�Ph�f �������������������U��h�jh�f �̙������t
�@��t]�����]�������U��Vh�jh�f 蛙��������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R��y���E�NP�у�4�M����y����^]ÍM��y�����^]��U��h�jh�f �,�������t
�@��t]��3�]��������U��h�jh�f ���������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á���H�F��  h�Tj8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��S�]V��F;�~ ��x�F�M��^�   []� ^3�[]� }jW�F9FuK��u�~��N�<��u�< ��tA����B�V��  h�Tj8��    QR�Ѓ���t�F�~�N�V��    �F9^|�_�F;Fu���������u����N�V�E���   F^[]� ��U��V��FW�};�~����y3�;Fu�m�����u_^]� �F;�~�N�T����H�;��F�M���F_�   ^]� ����U��E��x2�Q;�}+J�Q;�}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�c:��3����_�F�F^�����A    ��������̋Q�B���x;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�U�m8��3����_�F�F^��������������U���SV�uW���^S�}��68��3���F�F�O�N�W���V�E9G~|��I �O���F�U�9FuL��u�~��~��t���< ��tY����H���  h�Tj8��    RP�у���t0�~�}���V��M����E�F@�E;G|�_^�   [��]� _^3�[��]� U��V�u��x'�A;�} �U��x;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��x,�Q;�}%��x!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|����Ѕ�x);�}%N�q;�}�A�t���B�0;Q|�_�   ^]� _3�^]� ������U����E�Qj�E��ARP�M��E�U論����]� �����U����Q�Ej�E��A�MRPQ�M��E�U�ǖ����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q��T��t!�A��t�B�A�Q�P�A    �A    �̋�� U�@�T�HV3��q�q�P�r�r��T�p�p�p�P�H^������V���U�r����F3��F�T;�t�N;�t�H�F�N�H�V�V�F�F�T;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3���T;�t�F;�t�A�F�N�H�V�V�Et	V��7������^]� ������������U��V��W�~W�U�4��3����E��F�Ft	V�7����_��^]� ������U��V��������Et	V�7������^]� ���������������U�����PH�EPQ���  �у�]� �U�����P�B4VW�}j��h�  ���ЋMWQ���T  _^]� ��������������U��V���PXW�ҋ}P����������Et�_�   ^]� �M�UPWQR���A  _^]� �����������U��S�]VW��j �������8�  �}uI�~ uC����P���   j h�  ���Ѕ�u����QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ����  _^[]� ��������U��EP�A    �]Z����]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �y  ����   �M3�V�����8�  u4�]Q��P�w��Y������P�M�B4��jh�  ��_^�C�[��]� �MV�e����8�  u�E�M��RPQ����_^�   [��]� �MV�5����8�  t�MV�$����8��  ����P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P��,��3��؃��u�;�t����QH���  VS�Ѓ��E��M�;O�b  9w�Y  ����B�M���   Vh�  �҅�u!����P�M���   Vh�  �Ѕ��  ����Q�M�B4Vh�  ��;�t
V���������E��G������   ���   �Ћ]�E�;���   ;���   S�W���M���jQ�ˉu��uĉuȉủuЉu؉u��B=���U�E��ˉu��u�u�U�E��]��E�   �\L����tHtHt�u���E�   ��E�   ��E�   �����M�;�t�P����BX�M�Q����P������M܃�;�t�P���M�������M�������M��hX���]�U�E�MRSPQ���  _^[��]� ������   ���   �E�P�у�_^�   [��]� ��������������̸   � ��������� ������������̃��� ����������� �������������U�����H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ����Q0�F�M���   PQW�ҋF��^_]� U�����H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U�����H���  ]��������������U�����H���  ]��������������U�����P�EP�EP�EP�EPQ���   �у�]� �����U�����E�P�EP�E���\$�E�$PQ���   �у�]� �������������U�����P�EP�EP�EPQ���   �у�]� ��������̡���P���   Q�Ѓ�������������U�����P�EP�EP�EPQ���   �у�]� ���������U�����P�EP�EPQ���   �у�]� �������������U�����H�U�ApR�Ѓ�]� �����U�����P�EP�EPQ���  �у�]� �������������U�����P�EP�EPQ���  �у�]� �������������U�����P�EP�EPQ���  �у�]� �������������U�����P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P�t  ��R���E�P���ҡ���P�B<�M��Ћ}��t0j �M�QW���������u����B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4���� �E�py�E� � �E�0� �E��y�E�Р �E��y�E� � ǅx����yǅ|���`y�E�� �E�@� �E��� �E��y�E��y�E�Py�E�`� �E��� �E��y�E�� �E�P� �(���������B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u����H�A�UR�Ѓ�^3�[��]Ë���Q�B<W�M3��Ѕ��N  謭���E�����   �MQ�M���e������B�P�M�Q�ҡ���H�AWj��U�h�SR�Ѓ��M�Q�M��e���u�Wj��U�R�E�P��\���Q�_?�x����P��x���R�i����P�E�P�i����P���Ʈ���E���t�E� �� t�M������e����t��x��������e����t��\�������e����t�M̃���e����t����Q�J�E�P����у���t�M��ye���}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�x�������E$�M�UVP�Ej QRP�������������Q�J�EP�у���_^[��]���������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`L����������̋�`����������̋�` ����������̋�`����������̋�`D����������̋�`����������̋�`H����������̋�`����������̋�`,��U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E�9zj �u�u��u�i�  �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�  �� �E�_^[�E���]Ë�U��V��u�N3��  j V�v�vj �u�v�u��  �� ^]Ë�U���8S�}#  u�v{�M�3�@�   �e� �Eܢ{�8��M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E���  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����+���u�O  �MN��k�E�9H};H~���u	�M�]�u�} }̋EF�0�E�;_w;�v�  ��k�E�_^[�Ë�U��EV�u��n  ���   �F�`  ���   ��^]Ë�U���K  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�#  �u;��   u�  �N���   ^]��  ���   �	�H;�t���x u�^]�b  �N�H�ҋ�U����8��e� �M�3��M�E��E�E�E@�E�z�M��E�d�    �E�E�d�    �uQ�u�V  �ȋE�d�    ����;8�u���  ����Б�ԑy��ؑ-��ܑf����Ϟ�����������M����ٝË�U�������} t�*  ��]���������������̃��$�]-  �   ��ÍT$�-  R��<$�D$tQf�<$t��,  �   �u���=� �3-  �   �P��0-  �  �u,��� u%�|$ u���,  �"��� u�|$ u�%   �t����-V�   �=� ��,  �   �P���+  Z������̃=<� t-U�������$�,$�Ã=<� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̃=4� ��/  ���\$�D$%�  =�  u�<$f�$f��f���d$��/  � �~D$f(@Uf(�f(�fs�4f~�fTpUf��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�R,  ���D$��~D$f��f(�f��=�  |!=2  �fT0U�\�f�L$�D$����f�`UfV`UfTPUf�\$�D$Ë�Q��U�/  YË�U��V��������EtV�#��Y��^]� ��U��E��	Q��	P��/  ��Y�Y@]� jhX}��:  �E��uz�~:  ��u3��8  �  ��u�:  ���:  �P�@��k9  ���3  ��y�=  ���8  ��x �6  ��xj �Z1  Y��u����   �5  ��3�;�u[9=�~����}�9=��u�3  9}u�t5  ��  ��9  �E������   �   3�9}u�=���t�  ��j��uY�l  h  j�/  YY��;�����V�5���5,��P�Ѕ�tWV�  YY�P��N��V��  Y�������uW��  Y3�@�9  � jhx}�^9  ����]3�@�E��u9���   �e� ;�t��u.��U��tWVS�ЉE�}� ��   WVS�C����E����   WVS�.����E��u$��u WPS����Wj S������U��tWj S�Ѕ�t��u&WVS�������u!E�}� t��U��tWVS�ЉE��E������E���E��	PQ��;  YYËe��E�����3��8  Ë�U��}u�;  �u�M�U�����Y]� ��U��QSV�5PW�5(����5$��؉]��֋�;���   ��+��G��ruS��<  �؍GY;�sH�   ;�s���;�rP�u���-  YY��u�C;�r>P�u���-  YY��t/��P�4��P�(��u�=P�׉��V�ף$��E�3�_^[�Ë�Vjj �L-  YY��V�P�(��$���ujX^Ã& 3�^�jh�}�^7  ��-  �e� �u�����Y�E��E������	   �E��z7  ���-  Ë�U���u���������YH]��������U��WV�u�M�}�����;�v;���  ���   r�=<� tWV����;�^_u�>  ��   u������r)��$�`��Ǻ   ��r����$�t��$�p���$�������ԅ#ъ��F�G�F���G������r���$�`��I #ъ��F���G������r���$�`��#ъ���������r���$�`��I W�D�<�4�,�$����D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�`���p�x������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$����I �Ǻ   ��r��+��$� ��$�����4�\��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I ������ȇЇ؇����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�������$�8��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������̋T$�L$��ti3��D$��u���   r�=<� t�;  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$Ë�U��S�]���woVW�=�� u� :  j�J8  h�   �y)  YY��t���3�@Pj �5���P����u&j^9�tS�[<  Y��u����;  �0��;  �0��_^�S�:<  Y��;  �    3�[]Ë�U��} t-�uj �5���P��uV�;  ���PP�[;  Y�^]���U��<  ��U��V����U��<  �EtV����Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR��&  YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =RCC�t=MOC�t=csm�u*��  ���    ��  ��  ���    ~�  ���   3�]�jh�}�l1  �}�]��   �s��s�u��  ���   �e� ;utb���~;w|��  �ƋO�4��u��E�   �|� t�sh  S�O�t��   �e� ��u��+���YËe�e� �}�]�u��u���E������   ;ut�x  �s�1  Ë]�u���  ���    ~��  ���   Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�  3�A��  ���3��jh�}�K0  �M��t*�9csm�u"�A��t�@��t�e� P�q�(����E������Z0  �3�8E��Ëe��j  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�{  �*  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�^�������u
K�������E��E��E�;|�^[�E���j��G�/:  �  ���    t��  �e� ��  �M���  �]  �Mj j ���   �):  �j,hX~�	/  �ً}�u�]�e� �G��E��v�E�P����YY�E��  ���   �E��  ���   �E���
  ���   ��
  �M���   �e� 3�@�E�E��u�uS�uW��������E�e� �o�E������Ëe��
  ��   �u�}�~�   �O��O�^�e� �E�;Fsk��T;�~A;L;�F�L�QVj W�������e� �e� �u�E������E    �   �E��@.  ��E�맋}�u�E܉G��u������Y�
  �Mԉ��   �
  �MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v�j���Y��t�uV�%���YY�jh�~�m-  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w�z8  YY����   SV�i8  YY����   �G��M��QP�����YY���   �}�E�p�tH�28  YY����   SV�!8  YY����   �w�E�pV�)8  �����   ���t|��W�9Wu8��7  YY��taSV��7  YY��tT�w��W�E�p�_���YYPV��7  ���9�7  YY��t)SV�7  YY��t�w�7  Y��t�j X��@�E����  �E������E��3�@Ëe��i  3��@,  �jh�~��+  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS������FP�w����YYP�vS�����E������+  �3�@Ëe���
  ̋�U��} t�uSV�u�V������}  �uuV��u �G����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�����]Ë�U���V�u�>  ���   W�  ���    tG�  ���   �H  9t3�=MOC�t*=RCC�t#�u$�u �u�u�u�uV�b���������   �}� u�1
  �u�E�P�E�PV�u W�����M���;M�sg���E�S�x�;7|G;p�B���H�Q��t�z u-�Y��@u%�u$�u�u j �u�u�u�u�����u�E����E��M����E�;M�r�[_^�Ë�U���4�MS�]�CVW�E� =�   �I��I�M����|;�|�m	  �u�csm�9>��  �~� ��)  �F;�t=!�t="��  �~ �  �  ���    ��  �  ���   �u�  ���   jV�E�4  YY��u��  9>u&�~u �F;�t=!�t="�u�~ u��  �=  ���    ��   �+  ���   �   �u3����   ����Y��u\3�9~�G�Lh���������uF��;7|��  j�u�M���YY�EP�M��E�U�2  h�~�E�P�E̔U�3  �u�csm�9>��  �~��  �F;�t=!�t="���  �}� ��   �E�P�E�P�u��u W�g����M���;M���   �x�}�M��G��E�9��   ;O���   ��E�G��E��~r�F�@�X� �E��~#�v�P�u�E���������u�M��9E���M�E��}� ��.�u$�}��u �]��u��E��u�u�uV�u�����u�}���E��E����}�;E��P����}�} t
jV�����YY�}� ��   �%���=!���   �����   V�H���Y����   �H  �C  �>  ���   �3  �}$ �M���   Vu�u��u$������uj�V�u�u�X������v�g����]�{ v&�} ������u$�u �u�S�u�u�uV������ ��  ���    t�6  _^[�Ë�U��V�u���&1  ��U��^]� ��U��SVW�  ��   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�z������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������ 3�@_^[]�j �P�� P� ��V�5���$P����u�5(��P��V�5���(P��^á�����tP�50��P�Ѓ���������tP�,P�����#4  jh��$  h�U�4P�u�F\pW�f 3�G�~�~pƆ�   CƆK  C�Fh@�j�	5  Y�e� �vh�0P�E������>   j��4  Y�}��E�Fl��u�8��Fl�vl��4  Y�E������   �$  �3�G�uj��3  Y�j��3  YË�VW�P�5����������Ћ���uNh  j��  ��YY��t:V�5���5,��P�Ѕ�tj V�����YY�P�N���	V�H���Y3�W�8P_��^Ë�V��������uj�  Y��^�jh8�#  �u����   �F$��tP�����Y�F,��tP�����Y�F4��tP�����Y�F<��tP�����Y�F@��tP�����Y�FD��tP����Y�FH��tP����Y�F\=pWtP����Yj�{3  Y�e� �~h��tW�<P��u��@�tW�i���Y�E������W   j�B3  Y�E�   �~l��t#W��3  Y;=8�t��`�t�? uW�l4  Y�E������   V����Y��"  � �uj�2  YËuj�2  YË�U��=���tK�} u'V�5���5$P�օ�t�5���5�����ЉE^j �5���5,��P���u�x���������t	j P�(P]Ë�Wh�U�4P����u	�����3�_�V�5@Ph�UW��h�UW�$���h�UW�(���h�UW�,��փ=$� �5(P�0�t�=(� t�=,� t��u$�$P�(��,P�$����5,��0�� P��������   �5(�P�օ���   ��  �5$��5P���5(��$����5,��(����50��,��֣0���/  ��tc�=PhO��5$����У�����tDh  j�  ��YY��t0V�5���5,����Ѕ�tj V����YY�P�N��3�@��i���3�^_�jh`�   �����@x��t�e� ���3�@Ëe��E������V%  �   ������@|��t������jh��A   �54��P��t�e� ���3�@Ëe��E������}����hg��P�4������U���SQ�E���E��EU�u�M�m��;  VW��_^��]�MU���   u�   Q�w;  ]Y[�� ��U���(  �@��<��8��4��50��=,�f�X�f�L�f�(�f�$�f�% �f�-���P��E �D��E�H��E�T����������  �H��D��8�	 ��<�   �8��������<��������TP���j��:  Yj �PPh�U�LP�=�� uj�:  Yh	 ��HPP�DP�Ë�U��EV���F ��uc������F�Hl��Hh�N�;8�t�p��Hpu�1  ��F;h�t�F�p��Hpu�84  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P�R=  ��e�F�P� <  ��Yu��P�5=  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�p<  �M��E��M��H��EP��<  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�z=  @PV�V�(  ��^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M�������3�;�u"�%  j^�0��9  �}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�V%  j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]h�USV��<  ����ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F�X�_t�90uj�APQ�&  ���}� t�E��`p�3������3�PPPPP�i8  ̋�U���,�8�3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0��=  ����u�$  ��s8  ���m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q�;<  ����t� ��u�E�j P�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �Y���9}}�}�u;�u#�2#  j^�0�7  �}� t�E�`p����  9}v؋E��� 9Ew	��"  j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V�5  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� ��<  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �y<  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���W�<  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP��:  0�F�U�����;�u��|��drj jdRP�:  0��U�F����;�u��|��
rj j
RP�:  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u���w�ٍM�N�������u#��  j^�0�,4  �}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^�7  @PVS�!  �0�������} ~QV�^��6  @PVS�!  �E����   � � ������y&�߀} u9}|�}�}������Wj0S�*������}� t�E��`p�3�_^[�Ë�U���,�8�3ŉE��EVW�}j^V�M�Q�M�Q�p�0�8  ����u�  �0�3  ���lS�]��u�  �0��2  ���S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P��6  ����t� ��u�E�j VS���N�����[�M�_3�^�����Ë�U���,�8�3ŉE��EV�uWj_W�M�Q�M�Q�p�0��7  ����u��  �8�V2  ���   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW�16  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u��������u�E�jP�u���u�u������[�M�_3�^������Ë�U��E��et_��EtZ��fu�u �u�u�u�u�'�����]Ã�at��At�u �u�u�u�u�u������0�u �u�u�u�u�u�o�����u �u�u�u�u�u�o�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3���Б�P��Б����(r�_^Ë�Vh   h   3�V��7  ����t
VVVVV�f0  ^���������������̀zuf��\���������?�f�?f��^���٭^����,V�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����,V�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����$V���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-V��p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�6  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��@V�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��lV�����������\V�����   s��|V��dV�����������TV�����   v��tV�j
�XP�<�3�Ë�U���(3��E��E�9\�t�58��P��V��M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �E�DW�M��M�u�]���M��]�Q��]���Y����  �  � "   ��  �E�@W�M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �E�@W��E�8W�M�u��M�]���]���?  �U��E�8W�W����E�4W�ΉU��E�4W�?����E�DW�q�����tWItHIt9It ��t���  �E�,W��E�$W��E�DW�M��u��u����E�DW�c����E�   �������E���   �E�   �E�W�������������   �$�d��E�4W��E�8W��E�@W��E�W��E�W�t����E�W�h����E��V�\����E��V��E��V��E��V�M��u�M����M�]���]�M��]�Q�E�   ��Y��u��  � !   �E��^�Ð��ɮҮۮ��s���T�K����j
�XP�4�3�Ë�U��QQSV���  V�5 ��%;  �EYY�M�ظ�  #�QQ�$f;�uU�9  YY��~-��~��u#�ESQQ�$j�:8  ���tVS��:  �EYY�f�ES��Q���\$�E�$jj�A�$9  �]��E�Y�EY������DzVS�:  �E�YY�"�� u��E�S���\$�E�$jj�8  ��^[��jh��t  j��  Y�e� �u�N��t/�d��`��E��t9u,�H�JP����Y�v����Y�f �E������
   �c  Ë���j�  YËT$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U��VW3��u�Q�����Y��u'9h�vV�\P���  ;h�v��������uʋ�_^]Ë�U��VW3�j �u�u�_;  ������u'9h�vV�\P���  ;h�v��������uË�_^]Ë�U��VW3��u�u�;  ��YY��u,9Et'9h�vV�\P���  ;h�v��������u���_^]Ë�U��hXW�4P��thHWP�@P��t�u��]Ë�U���u�����Y�u�`P�j�  Y�j��  YË�V�������V��  V�[%  V�i  V�=  V�;  V������^Ë�U��V�u3����u���t�у�;ur�^]Ë�U��= U th U��=  Y��t
�u� UY�w���h(QhQ����YY��uTVWh�������Q�QY��;�s���t�Ѓ�;�r�=0� _^th0��=  Y��tj jj �0�3�]�j h��Z  j�  Y�e� 3�@9����   ����E����} ��   �5(��5P�֋؉]Ѕ�th�5$��֋��}ԉ]܉}؃��}�;�rK�t���9t�;�r>�7�֋��a�������5(��֋��5$���9]�u9E�t�]܉]ЉE؋��}ԋ]���E�,Q�}�8Qs�E� ��t�ЃE����E�<Q�}�@Qs�E�� ��t�ЃE����E������    �} u)���   j��  Y�u�����} tj�  Y��l  Ë�U��j j�u������]�jj j ������Ë�U����  �u�8  Yh�   ����̋�U���LV�E�P�tPj@j ^V����YY3�;�u����  ��   � ��5�;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5 ���@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9�}k�$�j@j �����YY��tQ�� ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9�|����3���~r�E�� ���t\���tW�M��	��tM��uP�pP��t=����������4� ��E�� ��E�� �Fh�  �FP�lP����   �F�E�G�E�;�|�3ۋ���5 �����t���t�N��q�F���uj�X�
�C�������P�hP�����tB��t>W�pP��t3%�   �>��u�N@�	��u�Nh�  �FP�lP��t,�F�
�N@�����C���h����5��dP3�_[^�Ã������VW� ����t6��   ;�s!�p�~� tV�xP���@   �N�;�r��7������' Y���� �|�_^Ã=,� u��  V�5�W3���u����   <=tGV��$  Y�t���u�jGW�������YY�=|���tˋ5�S�3V�$  �>=Y�Xt"jS����YY���t?VSP�%%  ����uG���> u��5������%� �' � �   3�Y[_^��5|�������%|� �����3�PPPPP��   ̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�49  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�O8  Y��t��M�E�F��M��E���,8  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9,�u�H  h  ���VS����|P�@��5��;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H�p��5t�3�����_^[�Ë�U���SV��P��3�;�u3��wf93t��f90u���f90u�W�=�PVVV+�V��@PSVV�E��׉E�;�t8P�;���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u�����Y�u�S��P�E��	S��P3�_^[�Ë�V��{��{W��;�s���t�Ѓ�;�r�_^Ë�V��{��{W��;�s���t�Ѓ�;�r�_^�j h   j ��P3Ʌ����������5����P�%�� ������h`�d�5    �D$�l$�l$+�SVW�8�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s358�W��E� �E�   �{���t�N�38� ����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t����/  �E���x@G�E��؃��u΀}� t$����t�N�38�����N�V�3:�����E�_^[��]��E�    �ɋM�9csm�u)�=�U t h�U�3  ����t�UjR��U���M�U�/  �E9Xth8�W�Ӌ��/  �E�M��H����t�N�38�����N�V�3:������E��H���/  �����9S�O���h8�W���1/  ������U��V����������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����8��e� �e� SW�N�@��  ��;�t��t	�У<��eV�E�P��P�u�3u���P3��P3���P3��E�P��P�E�3E�3�;�u�O�@����u��G  ����58��։5<�^_[�Ë�U��� �e� Wj3�Y�}��9Eu�*  �    �  ����x�MV�u��t��u�  �    �c  ����S�����E�;�w�M��u�E��u�E�B   �u�u�P�u���3  ������t�M�x�E��  ��E�Pj �1  YY��^_�Ë�U���uj �u�u�u�<�����]Ë�U��} u�r  �    ��  ���]��uj �5����P]���-  ��tj��-  Y�P�tjh  @j�  ��j����̋�U��3��M;Ő`t
@��r�3�]ËŔ`]Ë�U����  �8�3ŉE�SV�uWV������3�Y�����;��l  j�A  Y���  j�A  Y��u�= ���   ���   �6  h�ah  ���W��@  ������   h  ��VSf����P��  ��uh�aSV�@  ����t3�PPPPP�B  V�@  @Y��<v*V�v@  �El���+�j��h�a+�SP�?  ����u�h�a�  VW��>  ����u������VW��>  ����u�h  h@aW�h=  ���^SSSSS�y���j��hP��;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]���  YP�����PV��P�M�_^3�[�ú����j�@  Y��tj�@  Y��u�= �uh�   �%���h�   ����YYË�U��E�خ]�W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U�����U��E3�;�X�tA��-r�H��wjX]Ë�\�]�D���jY;��#���]��x�����u���Ã���e�����u�ēÃ�Ë�U��V������MQ�����Y�������0^]Ë�U��E�ܮ]Ë�U���5ܮ�P��t�u��Y��t3�@]�3�]ËA��u�bË�U��} W��t-V�u��  �pV�����YY�G��t�uVP�\  ���G^_]� ��V��~ t	�v�O���Y�f �F ^Ë�U��EV��f �b�F �0������^]� ��U��V�uW��;�t�����~ t�v���V�����F�G��_^]� �b�{�����U��V���b�h����EtV�����Y��^]� ��U��V�u��f �b�F �{�����^]� Pd�5    �D$+d$SVW�(��8�3�P�e��u��E������E�d�    Ë�U��� �EVWjY� b�}��E��E_�E�^��t� t�E� @��E�P�u��u��u���P�� ��U��3�@�} u3�]����������������U��WV�u�M�}�����;�v;���  ���   r�=<� tWV����;�^_u�|�����   u������r)��$����Ǻ   ��r����$���$� ���$�����@�d�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$����� ���(��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�<��I �Ǻ   ��r��+��$����$�����������F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I @�H�P�X�`�h�p����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�VW3����<�ԓu��Г�8h�  �0���lP��tF��$|�3�@_^Ã$�Г 3����S�xPV�ГW�>��t�~tW��W�����& Y�����|ܾГ_���t	�~uP�Ӄ����|�^[Ë�U��E�4�Г��P]�jh��[���3�G�}�3�9��u�>���j����h�   ����YY�u�4�Г9t���mj����Y��;�u�M����    3��Pj
�X   Y�]�9u+h�  W�lP��uW�M���Y�����    �]���>�W�2���Y�E������	   �E�������j
�)���YË�U��EV�4�Г�> uP�#���Y��uj�}���Y�6��P^]Ë�U��SV�50PW�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5<PW�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=Нth���   ;�t^9uZ���   ;�t9uP�x������   �X9  YY���   ;�t9uP�W������   ��8  YY���   �?������   �4���YY���   ;�tD9u@���   -�   P�������   ��   +�P� ������   +�P�������   ���������   =��t9��   uP��4  ���   辺��YY�~P�E   ���t�;�t9uP虺��Y9_�t�G;�t9uP肺��Y���Mu�V�s���Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu��`�tV�s���Y��^�3�_]�jh ������������p��Fpt"�~l t�����pl��uj �{���Y�������j�����Y�e� �58���lV�Y���YY�E��E������   �j�����Y�u��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�S���3��ȋ��~�~�~����~����@����F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �8�3ŉE�SW������P�v��P�   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R萷�����C����u�j �v�������vPW������Pjj �n:  3�S�v������WPW������PW�vS�!9  ��DS�v������WPW������Ph   �vS��8  ��$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�ѫ����jh ��
����:������p��Gpt�l t�wh��uj �����Y���"����j�0���Y�e� �wh�u�;5h�t6��tV�<P��u��@�tV����Y�h��Gh�5h��u�V�0P�E������   뎋u�j�����YË�U���S3�S�M������8����u�8�   ��P8]�tE�M��ap��<���u�8�   ��P�ۃ��u�E��@�8�   ��8]�t�E��`p���[�Ë�U��� �8�3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�p���   �E��0=�   r����  �t  ����  �h  ��P��P���V  �E�PW��P���7  h  �CVP賴��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�l����M��k�0�u������u��+�F��t)�>����E���l�D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C��t�Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����958��T�������M�_^3�[�Ȩ����jh@������M���-������}�������_h�u�q����E;C�W  h   �E���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�<P��u�Fh=@�tP����Y�^hS�=0P���Fp��   �p���   j����Y�e� �C�H��C�L��C�P�3��E��}f�LCf�E<�@��3��E�=  }�L��`�@��3��E�=   }��  ��h�@���5h��<P��u�h�=@�tP�2���Y�h�S���E������   �0j�'���Y��%���u ��@�tS�����Y������    ��e� �E�����Ã=,� uj��V���Y�,�   3�������U��SVWUj j h���u��n  ]_^[��]ËL$�A   �   t2�D$�H�3��ɦ��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    �8�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ�`��SQ�`��L$�K�C�kUQPXY]Y[� ��Ã%� ��U��W�}3�������ك��E���8t3�����_�Ë�U��E�T�]Ë�U���(  �8�3ŉE�S�]W���tS����Y������ jL������j P�������������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M�������������TPj ���PP������P�LP��u��u���tS����Y�M�_3�[�f����Ë�Vj� �Vj�������V�HPP�DP^Ë�U���5T��P��t]���u�u�u�u�u�����3�PPPPP�������Ë�U����u�M������E����   ~�E�Pj�u��1  ������   �M�H���}� t�M��ap��Ë�U��=̰ u�E�(��A��]�j �u����YY]Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS�<1  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�1  YY��t�Ej�E��]��E� Y��R���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�!/  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=̰ u�E�H���w�� ]�j �u�����YY]Ë�U���(�8�3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�;  �E�E�VP��0  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[蜡���Ë�U���(�8�3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P��:  �E�E�VP�5  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[���������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��UVW��t�}��u�����j^�0�(������3�E��u����+���@��tOu��u� ����j"Y�����3�_^]Ë�U��MS�YV�u3�;�u�j���j^�0��������   9Ev�U�;�~��@9Ew�>���j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W�v���@PWV������3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0�8�3ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f���>  �u܉C�E��E��C�E�P�uV�������$��u�M�_�s^��3�[������3�PPPPP�������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�I���YË�U��E�M%����#�V�u������t$��tj j �oG  YY��S���j^�0�������P�u��t	�KG  ���BG  YY3�^]Ë�S��QQ�����U�k�l$���   �8�3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�(  ��h��  ��x�����  �>YYt�=�� uV�    Y��u�6��  Y�M�_3�^�j�����]��[�3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�c  �EPSj �u��P�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�  Y����  �t�Etj�y  Y����x  ����   �E��   j�W  �EY�   #�tT=   t7=   t;�ub��M��������{L�H��M�����{,����2��M�����z������M�����z�p���p���������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�  �M��]�� �����������}�E����Q�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj�   Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}������ "   ]������� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3��ň�;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�S�������uV�,���Y�E�^�ËŌ��h��  �u(�  �u�����E ���Ë�U��=�� u(�u�E���\$���\$�E�$�uj�/�����$]������h��  �u� !   �\  �EYY]Ë�S��QQ�����U�k�l$���   �8�3ŉE��s �CP�s��������u#�e��P�CP�CP�s�C �sP�E�P�j������s�o������=�� u+��t'�s �C���\$���\$�C�$�sP�q�����$�P�����$��  �s �  �CYY�M�3��d�����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������&Q���EQQ�$������U�����  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-���]���t����-���]�������t
�-���]����t	�������؛�� t���]����jh`�����3�9<�tV�E@tH9��t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�� �e��U�E�������e��U�j��������SVW�T$�D$�L$URPQQhp�d�5    �8�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�r����   �C�����d�    ��_^[ËL$�A   �   t3�D$�H3��)���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�����3�3�3�3�3���U��SVWj Rh�Q�X  _^[]�U�l$RQ�t$������]� ��U��M��tj�3�X��;Es������    3�]��MV���uF3����wVj�5���P��u2�=� tV�	���Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u����Y]�V�u��u�u蔛��Y3��MW�0��uFV�uj �5����P����u^9�t@V����Y��t���v�V�z���Y�����    3�_^]��������PP����Y�����������PP����Y����ʋ�U��E������������]Ë�U��E�XV9Pt��k�u��;�r�k�M^;�s9Pt3�]��5���P�j h���1���3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC��������}؅�u����T  �������U�w\���]���Y�p��Q�Ã�t2��t!Ht�����    �^���빾�������������
�������E�   P�P�E�3��}���   9E�uj�D���9E�tP����Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,� X�M܋X X9M�}�M�k��W\�D�E����~�����E������   ��u�wdS�U�Y��]�}؃}� tj �K���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U��E���]�����������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h��h`�d�    P��SVW�8�1E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����u�M��s����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��QV�uV�RE  �E�FY��u������ 	   �N ����/  �@t������ "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�/C  �� ;�t�#C  ��@;�u�u�B  Y��uV�jB  Y�F  W��   �F�>�H��N+�I�N;�~WP�u�fA  ���E��M�� �F����y�M���t���t����������� �����@ tjSSQ�49  #����t%�F�M��3�GW�EP�u��@  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U��QSV�����`����G@� �E�t
� u�J�F����  �(�E� ��K�����E�>�u�'����8*u�ϰ?�u�����������8 u
�����M��^[�Ë�U���x  �8�3ŉE�S�]V�u3�W�u�}������������������������������������������������������������詨����u+�����    ����������� t
�������`p������
  �F@u^V�B  Y�����t���t�ȃ�������� �����A$u����t���t�ȃ������ �����@$��q���3�;��g����3ɉ��������������������������9
  G������9������&
  �B�<Xw����0m���3����Pmj��Y������;���	  �$�����������������������������������������������	  �� tJ��t6��t%HHt���u	  �������i	  �������]	  �������Q	  �������   �B	  �������6	  ��*u,���������[�������;��	  �������������	  ������k�
�ʍDЉ�������  ��������  ��*u&���������[�������;���  ��������  ������k�
�ʍDЉ������  ��ItU��htD��lt��w��  ������   �r  �?luG������   �������W  �������K  ������ �?  �<6u�4u�������� �  �������  <3u�2u�������������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������ ������P��P�  Y��������Yt"�����������������G������������������������������h  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@�������   ������������9������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  �������[���������  ;�u�ĝ������������ǅ����   �y  ��X��  HHty+��'���HH��  ��������  ������t0�C�Ph   ������P������P�?  ����tǅ����   ��C�������ǅ����   �������������/  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ���������P�����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�3���������T=  ���:��������� tf������f���������ǅ����   ��  ������@ǅ����
   �������� �  ��  ��S����  u��gucǅ����   �W9�����~�������������   ~=��������]  V�j���������Y��������t���������������
ǅ�����   ��5P���������C�������������P��������������������P������������WP�5����Ћ���������   t������ u������PW�5������YY������gu��u������PW�5�����YY�?-u������   G������W�
���ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �p���������Qƅ����0������ǅ����   �L�����   �R������� t��������@t�C���C����C���@t��3҉�������@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�7.  ��0���������ڃ�9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t��;�u�+��������(;�u����������������I�8 t@;�u�+����������������� �}  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+������������u'����~!������������� O�F����������t��ߋ�����������������P�������N���������Yt(������u��������ϰ0K������������t��ヽ���� ������tT��~P�������Pj�E�P������PK���E:  ����u ��������t�E�P�����������Y��u����������������������������Y������ |.������t%��������������ϰ K�H����������t��ヽ���� t����������������� Y���������������t������������3�������������� t
�������`p��������M�_^3�[��}���ÍI ������F����������U���$�8�3ŉE��ES�E��EVW�E��q����e� �=�� �E�u}hn��P�؅��  �=@PhnS�ׅ���   �5PP��h�mS�����P��h�mS�����P��h�mS�����P�֣����th�mS��P�֣������M�5P;�tG9��t?P���5�����֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3���;E�t)P�օ�t"�ЉE��t���;E�tP�օ�t�u��ЉE��5���օ�t�u�u��u��u����3��M�_^3�[�a|���Ë�U��V�uW��t�}��u�����j^�0�)�����_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f��y���j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�>���j^�0�������݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f�����j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u�n���j^�0�������_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f��.���j"Y���뼋�U��M��x��~��u��]á���]�������    �S������]Ë�U��E��t���8��  uP�����Y]Ë�U��V�u���c  �v�܅���v�ԅ���v�̅���v�ą���v輅���v贅���6譅���v 襅���v$蝅���v(蕅���v,荅���v0腅���v4�}����v�u����v8�m����v<�e�����@�v@�Z����vD�R����vH�J����vL�B����vP�:����vT�2����vX�*����v\�"����v`�����vd�����vh�
����vl�����vp������vt�����vx�����v|������@���   �Ԅ�����   �Ʉ�����   辄�����   賄�����   訄�����   蝄�����   蒄�����   臄�����   �|������   �q������   �f������   �[������   �P������   �E������   �:������   �/�����@���   �!������   �������   �������   � ������   ��������   �������   �߃�����   �ԃ�����   �Ƀ�����   较�����   賃�����   訃�����   蝃����   蒃����  臃����  �|�����@��  �n�����  �c�����  �X�����  �M�����  �B�����   �7�����$  �,�����(  �!�����,  ������0  ������4  � �����8  �������<  ������@  �߂����D  �Ԃ����H  �ɂ����@��L  軂����P  谂����T  襂����X  蚂����\  菂����`  脂����^]Ë�U��V�u��tY�;НtP�a���Y�F;ԝtP�O���Y�F;؝tP�=���Y�F0; �tP�+���Y�v4;5�tV����Y^]Ë�U��V�u����   �F;ܝtP����Y�F;��tP����Y�F;�tP�ρ��Y�F;�tP轁��Y�F;�tP諁��Y�F ;�tP虁��Y�F$;��tP臁��Y�F8;�tP�u���Y�F<;�tP�c���Y�F@;�tP�Q���Y�FD;�tP�?���Y�FH;�tP�-���Y�vL;5�tV����Y^]Ë�U����8�3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5�P3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w�X0  ��;�t� ��  �P����Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5�PSSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�/  ��;�th���  ���P���Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$��P�E�W�:���Y�u��1����E�Y�e�_^[�M�3��}s���Ë�U����u�M������u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap��Ë�U��QQ�8�3ŉE�S3�VW�]�9]u�E� �@�E�5�P3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w�\.  ��;�t� ��  �P��}��Y;�t	� ��  ���؅�t��?Pj S�8}����WS�u�uj�u�օ�t�uPS�u��P�E�S�����E�Y�e�_^[�M�3��Pr���Ë�U����u�M��ԑ���u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U���S�u�M�蓑���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�6����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M��ܐ���E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���8�8�3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=8�O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�4���+8�;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�58�N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��<��A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �<�;0���   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�D�0�3�@�   D��e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+<���M���Ɂ�   �ً@�]���@u�M̋U�Y��
�� u�M̉�M�_3�[�k���Ë�U���8�8�3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=P�O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�L���+P�;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5P�N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��T��A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �T�;H���   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�\�H�3�@�   \��e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+T���M���Ɂ�   �ًX�]���@u�M̋U�Y��
�� u�M̉�M�_3�[�kf���Ë�U���|�8�3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u袭���    �����3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$���Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  ����`�E�;���  }�عP��E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^��_���ÍI �2}��+?�� ����U���t�8�3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uh�v�S3�PPPPP�L���3�f9U�t��   �u9Uu-h�v�;�u"9Uuh�v�CjP��������u��C�h�v�CjP� �������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع���`�ۉE�f�U�u�}�M���  ��y�P���`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��V���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95<���  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��QQ�EV�u�E��EWV�E��W  ���Y;�u����� 	   �ǋ��J�u�M�Q�u�P��P�E�;�u�P��t	P����Y�ϋ����� ������D0� ��E��U�_^��jh���j�������]܉]��E���u覘���  苘��� 	   �Ë��   ��x;�r�~����  �c���� 	   ������ы����<� ���������L1��t�P��  Y�e� ��D0t�u�u�u�u��������E܉U������� 	   �	����  �]܉]��E������   �E܋U��܎����u�  YË�U���  �  �8�3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u蔗���8�z����    �׫������  ������S�� �������L8$�����$�����?�����t��u'�M����u�6����  �����    �x����  �D8 tjj j V������V�>  Y����  ��D���  ��i���@l3�9H�� �����P��4����P3�;��`  ;�t8�?����P  ��P��4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P����Y��t:��4���+�M3�@;���  j��D���SP�  �������  C��@����jS��D���P�  ������n  3�PPj�M�Qj��D���QP�� ���C��@�����P�����=  j ��,���PV�E�P��$���� �4��P���
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4��P����  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����+  Yf;�D����I  ��8�������� t)jXP��D�����  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4��P���C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4��P���i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  ��P��;���   j ��(���P��+�P��5����P��$���� �4��P��t�(���;����P��D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48��P��t��(�����D��� ��8�����P��D�����8��� ul��D��� t-j^9�D���u�<���� 	   �D����0�?��D����H���Y�1��$���� �D@t��4����8u3��$������    �����  ������8���+�0���[�M�_3�^�JI����jh��胇���]���u�Ȑ���  譐��� 	   ����   ��x;�r衐���  膐��� 	   �����ҋ����<� ��������D0��t�S��  Y�e� ��D0t�u�uS�n������E���,���� 	   �4����  �M���E������   �E�����Ë]S�?  YË�U���аh   �|��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u蟏��� 	   3�]Å�x;�r脏��� 	   �����ދȃ����� ����D��@]ø`�á �Vj^��u�   �;�}�ƣ �jP�{��YY����ujV�5 ��{��YY����ujX^�3ҹ`������� �����|�j�^3ҹp�W������ �����������t;�t��u�1�� B��О|�_3�^���
  �=�� t�  �5��R��YË�U��V�u�`�;�r"����w��+�����Q�v����N �  Y�
�� V��P^]Ë�U��E��}��P�I����E�H �  Y]ËE�� P��P]Ë�U��E�`�;�r=��w�`���+�����P�'���Y]Ã� P��P]Ë�U��M�E��}�`�����Q�����Y]Ã� P��P]Ë�U��E��u蕍���    �������]Ë@]á8���3�9԰����Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v�+���j^�0艡�����V�u�M��%e���E�9X��   f�E��   f;�v6;�t;�vWSV�	P���������� *   �Ռ��� 8]�t�M��ap�_^[��;�t&;�w 赌��j"^�0����8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p��P;�t9]�j����M;�t����P��z�P���;��s���;��k���WSV�>O�����[�����U��j �u�u�u�u������]����������Q�L$+ȃ����Y�  Q�L$+ȃ����Y�  ����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����ES3�VW�E�N@  ��X�X9]�E  �]����}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�K3�;�r��s3�B�ىH��t
�M�A�M�H�M�M�E�} �X�H�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[�Ë�U��MS3�VW;�|[;�sS��������<� �����D0t6�<0�t0�= �u+�tItIuSj��Sj��Sj���P���3���ڈ��� 	   ��������_^[]Ë�U��E���u�ƈ���  諈��� 	   ���]Å�x;�r袈���  臈��� 	   �����Ջ����� ������Dt͋]�jh �����}����������4� ��E�   3�9^u5j
�@���Y�]�9^uh�  �FP�lP��u�]��F�E������0   9]�t���������� ��D8P��P�E���~���3ۋ}j
����YË�U��E�ȃ����� ����DP��P]Ë�U��Q�=���u��  ������u���  ��j �M�Qj�MQP��P��t�f�E�Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��._���E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p��P���E�u�M;��   r 8^t���   8]��f����M��ap��Z�������� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p��P���:���뺋�U��j �u�u�u�������]������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��jh ��|��3ۉ]�j�����Y�]�j_�}�;= �}T����9�tE���@�tP��  Y���t�E��|(������ P�xP���4��I��Y����G��E������	   �E��h|���j蝋��YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�~���YP�O�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV����P�A  Y��Y��3�^]�jh@��]{��3��}�}�j詋��Y�}�3��u�;5 ���   ����98t^� �@�tVPV����YY3�B�U������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u���4�V�#���YY��E������   �}�E�t�E���z���j����Y�j����Y������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� 3�PPjPjh   @h�v��P���á�����t���tP��PË�U��V�uW�����u�?����    蜗����D�F�t8V�����V���N  V�p���P�~  ����y�����F��tP�&G���f Y�f ��_^]�jhh��y���M��3��u������u�ł���    �"��������F@t�f �E��y���V����Y�e� V�<���Y�E��E������   �ԋuV�e���Y�jh���)y���]���u�[���� 	   ����   ��x;�r�<���� 	   虖���ڋ����<� ��������D��t�S����Y�e� ��Dt1S�0���YP��P��u�P�E���e� �}� t�����M��Ł��� 	   �M���E������   �E��x��Ë]S�����Y�������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV�Y���Y���tP� ���u	���   u��u�@Dtj�.���j���%���YY;�tV����YP��P��u
�P���3�V�u��������� �����Y�D0 ��tW�Ā��Y����3�_^]�jh���Gw���]���u茀���  �q���� 	   ����   ��x;�r�e����  �J���� 	   觔���ҋ����<� ��������D0��t�S����Y�e� ��D0tS�����Y�E������� 	   �M���E������   �E���v��Ë]S����YË�U��V�u�F��t�t�v��C���f����3�Y��F�F^]��% P�������̍M������T$�B�J�3���7����{�4��������������̍M��	���M��P����T$�B�J�3��7����{�W4������̋E�P�^��YËT$�B�J�3��7���|�,4�����������̋E����   �e���M�����ËT$�B�J�3��O7���<|��3�������������̍M������M�������p����e���M��=����M��E����M�������@���������T����7���EP��]��YÍM��4���M��\����M��T����T$�B��|���3��6���`|�X3��������h`Rjh��E�P�{`����ËT$�B�J�3��6����|�3�������������̍M�������M�������M�������M�� X���T$�B�J�3��86���0}��2���T$�B�J�3��6���0~�2������������h�G�=��Y����̃=̣ uK�ģ��t����Q<P�B�Ѓ��ģ    �У��tV��� ���V�\�����У    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �� �� � "� 4� D� P� `� l� x� �� �� �� �� ʃ ڃ � � � ,� H� f� z� �� �� �� �� ΄ �� � � .� D� ^� t� �� �� �� ą ԅ � � � � 2� D� \� t� �� �� �� �� �� Ɔ ֆ � �� �  � 2� B� R� `� n�         �G        e��������5        �A�6                        failed to register EdgeSweep!        �f@-DT�!	@              �?objCopy �D�JW�?0x� P �� �� �� �� �� Н �  � �� � P� @� `� �  � �� �� �� �� �� �� �� � �� �� �� �� �� P� p� �   sweep_profile   edgeSpline  copy    _instance   ..\..\..\..\C4D 9.6\plugins\dev_complete\edgeSweep\source\tool\edgesweep.cpp    Oedgesweep  es.tif  EdgeSweep   n:\maxon\cinema4dr12demo\resource\_api\c4d_general.h    %s     n:\maxon\cinema4dr12demo\resource\_api\c4d_resource.cpp #   M_EDITOR    ����MbP?�x�� 0�  y�� n:\maxon\cinema4dr12demo\resource\_api\c4d_baseobject.cpp   Ly@� res     ������n:\maxon\cinema4dr12demo\resource\_api\c4d_file.cpp     �������      �?n:\maxon\cinema4dr12demo\resource\_api\c4d_libs\lib_ngon.cpp    n:\maxon\cinema4dr12demo\resource\_api\c4d_basebitmap.cpp   n:\maxon\cinema4dr12demo\resource\_api\c4d_pmain.cpp    `ypln:\maxon\cinema4dr12demo\resource\_api\c4d_gv\ge_mtools.cpp �y�l�yPl<z m(~                  �?      �?3      3            �      0C       �       ��              �z�    ���z����bad exception   K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    8���e+000                      ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �                  �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �      r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            0`   �_	   �_
   8_   �^   �^   8^   �]   p]    ]   �\   @\   �[   �[   �Z    �Z!   �Xx   pXy   TXz   8X�   0X�   XM i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     L{����Unknown exception   csm�               �        H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh     Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        �k�k�k�ktkhk\kTkLk@k4k1k,k$k kkkkkkk�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�j�jtjhj`jTj<j0jj�i�i�i�i|iXi<ii�h�h�h�h�h�h�hdh\hPh@h$hh�g�g�g`gDg g�f�f�f�f1ktfXfDf$ff( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx          GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L                                                                                                                                                                                                                                                                                       ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#QNAN  1#INF   1#IND   1#SNAN  C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           8�`{              �w�w�w     �       ����    @   �w�        ����    @   �w           �w�w               xx�w�w    0�       ����    @   �w            L�Dx           Txhxx�w�w    L�       ����    @   Dx           �x�x    d�        ����    @   �x            ���x           �x�x    ��        ����    @   �x            ��y           $y0y�x    ��       ����    @   y            ��w            ��ty           �y�y    ��        ����    @   ty            ؐ�y           �y�y    ؐ        ����    @   �y            ��z           z z�x    ��       ����    @   z            �Pz           `zhz    �        ����    @   Pz            `��z           �z�z    `�        ����    @   �z            ���z           �z�z{    ��       ����    @   �z��        ����    @   4{           D{{                ��4{�z �{ `� �� p� �E �E F YF �F )G pG �G                     �����E"�   �{                       �����E    �E"�   �{                       ����F"�   |                       ����@F"�   4|                       "�   �|                       �����F    �F�����F   �F   �F   �F   �F   �F   �F   �F   �F   �F����G"�   �|                       ����PG    XG   `G   hG"�   }                           ����    ����    ����    	�    ����    ����    ����i�z�    ����    ����    ����    ̄    ����    ����    ����    D�    ������    ����    �������@           ӌ����    ����                  �}"�   ~   ~                   ����    ����    ����    �    {�������    ����    �������    ����    ����    ��������    ��    �~   �~�~    ��    ����       ��    ��    ����       ������    ����    ����    ������    ������    ����    ����    f�����    r�����    ����    ��������    ����    ����    ����כۛ    ����    ����    ����    �    ����    ����    ����    Ŵ    ����    ����    ����    R�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    T�    ����    ����    ��������    ����    ����    ����    $�    ����    ����    ��������    ����    ����    ����    j-    ����    ����    ����    :5    ����    ����    ����    t=    ����    ����    ����    �?    ����    ����    ����    hA        4A����    ����    ����    �B    ����    ����    ����    �C    ����    ����    ����    fE�         ��  P                     �� �� � "� 4� D� P� `� l� x� �� �� �� �� ʃ ڃ � � � ,� H� f� z� �� �� �� �� ΄ �� � � .� D� ^� t� �� �� �� ą ԅ � � � � 2� D� \� t� �� �� �� �� �� Ɔ ֆ � �� �  � 2� B� R� `� n�     RtlUnwind �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer �HeapAlloc GetLastError  �HeapFree  �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  EGetProcAddress  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent IsProcessorFeaturePresent �Sleep ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �HeapSize  %WriteFile GetModuleFileNameW  �RaiseException  9LeaveCriticalSection  � EnterCriticalSection  rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage �HeapReAlloc ?LoadLibraryW  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  $WriteConsoleW � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll      �=�L              �� �� �� `b ԇ   edgesweep_R11.cdl c4d_main                                    �U    .?AVNodeData@@  �U    .?AVBaseData@@  �U    .?AVObjectData@@    �U    .?AVEdgeSweep@@ �U    .?AVGeSortAndSearch@@   �U    .?AVNeighbor@@  �U    .?AVDisjointNgonMesh@@  �U    .?AVGeToolNode2D@@  �U    .?AVGeToolDynArray@@    �U    .?AVGeToolDynArraySort@@    �U    .?AVGeToolList2D@@  N�@���Du�  s�          sqrt            �U    .?AVtype_info@@         �U    .?AVbad_exception@std@@ �U    .?AVexception@std@@ ��������            ��������������������        ?              �����
                                                                                                  	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                           C       �e�e�e�e|exetelede\ePeDe<e0e,e(e$e eeeeeeee e�d�d�d�de�d�d�d�d�d�d�d�d�d�dpddd	         \dTdLdDd<d4d,ddd�c�c�c�c�c�c�c�c�c�c�cxcpchc`cXcPc@c,c cc�cc�b�b�b�b�b�b�b�b|bTb@b                                                                                           �            �            �            �            �                              Н        (o�s0u��`�                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     @��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��     �            ����            �&         @W   DW   4W   8W    f   �e!   �e   ,W   $W   W   �e   �e   �V   �V    �V   W   W   �e   �V   �e   �e   �e   �e   �e"   �e#   �e$   �e%   �e&   �e      �      ���������              �       �D        � 0                 Dm4m.   .   ȝİİİİİİİİİ̝ȰȰȰȰȰȰȰН(o*q,q   ���5      @   �  �   ����              �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                                                                               �                 0  �              	  H   X� Z  �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel>
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPAD   �   00A0V0e00�0�0�0#1�1�1�12$2T2q2�2�2�2�2373M3a3r3}3�3�3�34-4H4u4�4�4�45T5j5�5�5�5�5�5�56&6A6G6M6Y6p6�6�6�6�67(7�7�7�78)8x8�8�8�89b9�9�9�9:�;�;4<T<�<=$=<=T=j=�=�=>,>?>P>w>�>�>�>�>??.?R?j??�?�?�?�?      �   0�0�0�011)1H1o1�1�1'2A263�3�3�3	4$4E4e4�4�5n6�6�7�7�7�7�78-8P8f8�8�8�8�8�89J9�9�9�9:.:Q:g:�:�:�:�:7;\;|;�;E<a<u<�<�<�<�<�<=*=o=�=�=�=�=�=>h>�>�>�>?>?U?c?}?�?�?�?   0  �   V0d0u0|0�0�0�0�0�01121c1u1�1�1�1�1�12212g2t2�2�2�2�23D3a3�3�3�34$4T4�4�4�45$5D5d5�5�5�5�5�56$6A6Q6d6�6�6�6�6!717D7�7�7�7�78!818A8T8t8�8�8�8�89?9d9�9�9�9�9�9:4:_:�:�:�:;*;T;t;�;�;�;�;<4<T<t<�<�<�<7=t=�=�=4>t>�>�>�>!?A?T?�?�?�?�?�?   @    0$0D0d0�0�0�01$1A1`1�1�1�1�1242t2�2�2�2�233&3T3t3�3�3�3�3 444D4d4�4�4�4�4-5;5N5c5�5�5�5�5�5�56"6D6l6�6�6�6�6�6$7<7e7~7�7�7�7�7�7848L8u8�8�8�8�8�899D9m9�9�9�9�9�9$:M:f:�:�:�:�:;$;D;o;�;�;�;�;<4<Q<d<�<�<�<�<=4=T=t=�=�=�=�=>4>Q>a>t>�>�>�>�>?$?9?K?T?e?{?�?�?�?�?�?   P  H  A0H0�0�0�01)1T1]1j1�1�1�1�1�1�1�1�12&2E2W2r2�2�2�2�2�233'393K3]3o3x3�3�3�3�3�34&484A4_4�4�4�4�4�455575I5[5m55�5�5�5�5�56$666H6Q6o6�6�6�6�6�6�67.7D7`7q7�7�7�7�7�7�7�788(8F8d8v8�8�8�8�8�8�8909F9b9t9�9�9�9�9�9 ::$:-:K:l:�:�:�:�:�:;!;�;�;�;�;�;�;�;<!<*<=<�<�<�<�<�<==D=a=�=�=�=�=>]>>�>�>�>�>�>?/?f?x?   `  �   0)0K0�0�0�1�12E2�2�2�2E3�3�3�34U4�4�4/5u5�5�5"6U6�6�627e7�7�7%8U8�8�8959�9�9:U:�:�:�: ;4;D;e;�;�;5<r<�<=E=�=�=	>1>Y>c>�>�>�>�>
?5?Y?�?�?�? p  �   0u0�0�01-1V11�1�1#2H2g2�2�2�213t3�3�3�3444a4�4�4�4�45A5d5�5�5�56^6�6�6�67$7D7t7�7�7�78!8D8t8�8�8�89D9d9�9�9�9�9:$:A:q:�:�:;d;�;�;�;�;<D<q<�<�<�<=1=Q=q=�=�=>$>T>�>�>�>?D?�?�?�?   �  �   !0A0a0�0�0�011141]1�1�1
242T2z2�2�273�3'4a4u4�4�4�45-5c5�5�5�5646T6�6�6P7�7�7�7�7$8Y8�8�8�8�89"9C9d9�9�9�9:!:D:d:�:�:;$;Q;q;�;�;�;<$<t<�<�<=$=D=�=�=�=�=1>N>x>�>�>�>?+?<?\?v?�?�?�?�? �  �   020o0�0�0�0�0+1>1a1{1�1�1�1�2�2�2�2<3D3i3�3�5o8�8�8�8 909g9�9�9t;x;|;�;�;�;�;<!<1<D<�<�<�<�<�<=$=L=�>�>�>;?�?�?�?�?�?�?�?�?�?�?   �  �   0000"0)000o1�1�1�12!2�2�2	3%3�3�3	4%4�4�4�4�45$5D5e5�5�5|6�6�6!7�7�7�7�78$818_8�8�8�8�899A9T9�9�9�9�9:":A:d:�:�:�:;4;Q;q;�;�;�;<4<a<�<�<�<�<1=Q=t=�=�=�=�=>4>T>t>�>�>�>�>?$?D?�?�?�?   �  �   \0�0�01a1�1�12�2�2�2Q3n3�3�3434�4�4515T5�5C6l6�67<7d7�7848�8�8�8[9�9�9Q:w:�:�:Q;w;�;<<�<�<=~=�=�=.>N>c>�>?|?�?   �  �   040Q0a0t0�0�0�0 1$1T1t1�1�1�1242Q2t2�2�23 3B3~3�3�3�344Q4q4�4�4�4�4�5�5�5�5�5�5646Q6d6�6�6�6747T7t7�7�7�7�78R8�8�8�8"9P9~9�97:N:{:�:�:;;�;	<<�<#>->7>A>K>U>_>t>�>�>�>??�?�? �  �   010T0t0�0�0�0�01D1d1�1�1�1�12;2a2�2"3a3�3�3�3�34$4T4f4�4�4�4�4$5D5a5�5�5�5�546�6�6747T7t7�7�7�7�78D8T8�8�8�8�8!9D9q9�9�9�9:A:d:�:�:�:;1;Q;q;�;�;�;�;<1<Q<q<�<�<�<�<=1=B=d=u=�=�=�=�=�=�=>!>2>T>t>�>�>�>�>�>? ?D?d?|?�?�?�?�?�?�? �  ,  00/0@0s0�0�0�0�0�0�01141T1t1�1�1�1�1�12D2d2�2�2�2�2313D3t3�3�3�3�34$4A4Q4a4t4�4�4�4�4545T5t5�5�5�5�560686L6�6�6�6717U7�7�7�7�7848T8t8�8�8�8�8919A9T9�9�9�9�9�9�9�9:3:A:P:q:�:�:�:�:;;!;1;D;d;;�;�;�;�;�;<$<D<d<�<�<�<�<=7=P=a=}=�=�=�=�=>>D>d>�>�>�>�>??/?>?N?`?�?�?�?�?�?�?   �  �   0(0N0e0|0�0�0�0�0�0�0121F1U1e1v1�1�122!242T2t2�2�2�2�2343T3t3�3�3�3�3444T4t4�4�4�4�45<5d5�5�5�5�5646T6t6�6�6�6�6747T7t7�7�7�7�7848T8t8�8�8�8�89$9D9d9�9�9�9�9�9�9:$:F:Z:j:�:�:�:�:�:;@;U;�;�;�;�;�;$<A<d<�<�<�<=    h   �01-1e1�1�152u2�2�2"3U3�3�34E4�4�4525b5�5�5�556u6�67U7�7�78e8�8%9;);�;.>�>�>�>�>�>�?�?�?�?   �   X0f0�0�0X1`1�1�1�1�13333A3�3�3�3�3�4�45$5A5T5�5�5�5�5646T6�6�6�6�6$7D7d7�7�788(8d8�8�8�89!9D9d9�9�9�9�9!:�:�:�:$;A;T;(=:=M=p=(?a?t?�?�?�? 0 �   !010S0t0�0�0�0171E1T1�1�1�1�1�1$2T283l3�3�3;4C5V5f566&6�6�6�6�7�7�7�7�7848T8t8�8�8�8�8�8�89$9D9d9�9�9�9�9:!:D:t:�:�:�:�:;4;T;t;�;�;�;�;<4<Q<o<�<�<�<�<=?=a=�=�=�=�=�=!>4>T>q>�>�>�>�>?5?r?�?�? @ �   u0�0�0E1�1�12b2�2�2%3e3�3�3%4�4�4�4b5�5�5�526b6�6�687h7|7�7�7�78U8�8�859�9�9%:u:�:;R;�;�;<b<�<%=b=�=%>b>�>�>E?�?�?   P x   50�0�0H1�1E2�2�23E3�3�324u4�45e5�5�5E6�6�6E7�7�7818]8�8�8%9e9�9:U:�:;U;�;<E<�<�<=U=�=�=5>�>�>?@?�?�?�?   ` x   \0�0�0<1�1�1@2F2t2�2�2�2�2�2�2"343N3d3h3l3p3t3x3�3�3�3D4t4�4�4�5�5�8}9�9�: ;�;�;�;�;�;<-<}<�<4=T=>$>�>v?�?�?   p �   000[0j1�1|2�2�3�3�3�344a4�4�4�4545d5�5�5(6}6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777X7u7�7�7�7�8�8%:�:�:�:b=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>>>#>�>�>�>�>�>?.?�?   � �   
0#0�0�0�0�0�051m1r1|1�1�1�1�12F2L2R2g2�2�2�2 3M3�3�3�384=4F4U4x4}4�4�45L5d5k5s5x5|5�5�5�5�5�5�5�5 66666Z6`6d6h6l6�6�6�6�6777-7W7�7�7�7�7�7�7�7�7�7�7�7 888�8�89!909�9�9�9�9�9�:�;�<�<�> �   	083h3r3}3�5�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6777%7G7\7�7�7�7�7�7�78,8R8�8�8�81999�9�9�9�9�9�9�9�9�9�9�9�9::::&:,:3:9:A:H:M:U:^:j:o:t:z:~:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;0;6;N;j;�;�;�;�;�;�;X<^<d<j<p<v<}<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<	===#=)=/=E=L=|=�=�=�= � �   Z0�0�0V67�8�8�8)9�98:�:k;l<|<�<�<�<�<�<�<�<�<�<�<^=�=�=�=>>>&>N>W>`>v>�>�>�>�>�>�>�>�>�>???d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?   � �   0�0�0�0�1�1�1�1�1�1,252A2]2c2l2s2�2
33%30353G3Q3V3r3|3�3�3�3�3�3�3�3�3*444Z4a4{4�4�4,5R5X5�5�5�5�5*646_6w6�6�6�6�6)7L7R7g7�7�7�7�7�78I8T8^8o8z8::K:S:Y:^:d:�:�:�:;f;r;�;�;�;�;�;�;�;�;�;<<r<L=T=l=�=�=b?�?�?�?�?�?�?�?�?   � �   �0�0101C1U1�1�1�1�1�1�1�1)262K2|2�2�23:3
5&5I5\5�5�5�5�5;6�6�6�6�6$7W7�7�7�7�7888898_8}8�8�8�8�8�8�8�8�8�8�8�8�8�8b9m9�9�9�9�9�9�9�9: :$:(:,:0:4:8:<:�:�:�:�:�:�:�:�:;";0;6;Y;`;y;�;�;�;�;�;<g<�<�<�<2=z=�=�>�>7?Q?b?�? � �   )0f0}0�1�182E2O2]2f2p2�2�2�2�2�2�23J33�344h4�4�4k5w5�5�5�5�5�5�5�566"6+606?6f6�6�6�6!7-7�7�7�7�7&8889"9/9m9t9�9�9::R;�;(<)? � p   51)24�5 66,646�6�78D8�8�8#;5;G;m;z;�;�;�;<=q=w=�=�=�=>8>P>j>o>t>y>�>�>�>�>??L?Q?X?]?d?i?w?�?�?�? � H   o011/1M1a1g1;3B3N4�45*5�5�5�59�9=;�;�;�;�=�?�?�?�?�?�?�?�?�?   x   0%0+0;0@0Q0Y0_0i0o0y00�0�0�0�0�0�0�0�01/11383>377%777I7o7�7�7�7�7�7�7�7�78#858G8`8�8B9:�:�:H;�<:=.>6>�>�?  `   `0f0111�1�12�23�3845�5�5X6^6l677Y7�7�:�:�= >>>>>>>> >$>(>5>�>?/?L?�?�?     $   �9I<V<o<�<�<�<�=�=�>�>�?�?   0 �   0�1`203a3w3�3�3t4�4�4L5�5�5�5�566!6-6=6D6S6_6l6�6�6�6�6�6�6(777@7d7�7�7�7�8�8<<2<R<�<�<�<=/=\=g=�=�=�=�=�=�>�>N?o?x?�?�?�?�?   @ \   �0�0�0�0:1�1�1�1�1�1Z2�2�23N3X3(4e4o4�4�4�4
5�5�56-6k6777;7�7�7�7�7�7�7�7�78   P �   1111 1$10141�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2`3d3h3l3p3�3�3�4�4555555 5�5�5�5�5�5�5�5�5 ` �   �0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1 222�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0= p D  |7�7�7�7�7�7�7�7�7�7�7 88888,8<8@8P8T8X8\8`8h8�8�8�8�8�8�8�8�8�8�8�899 9$9(909H9X9\9l9p9�9�9�9�9�9�9�9�9�9�9�9 :::: :8:H:L:\:`:h:�:�:�:�:�:�:�:�:�:�:�:�:�:;;0;@;D;X;\;�;�;�;�;�;<<8<D<h<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==$=,=8=p=�=�=�=�=�=�=�=�=>,>8>@>p>x>|>�>�>�>�>�>�>�>�>�>�>�>?(?4?P?\?t?x?�?�?�?�?�?   � ,   080X0t0x0�0�0�0�0�0181X1d1�1�1�1   � l   0000L0d0�0�0�0�0�01`1�1�1�1�1�1�1�1�1�1�1�1�1�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6�6�6�6�6�67(7,7074787h;�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>`>h>                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          